* Equivalent circuit model for TCM1-43X+_1.ckt
.SUBCKT TCM1-43X+_1 po1 po2 po3
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Vsp2 po2 p2 0
Vsr2 p2 pr2 0
Rp2 pr2 0 50
Ru2 u2 0 50
Fr2 u2 0 Vsr2 -1
Fu2 u2 0 Vsp2 -1
Ry2 y2 0 1
Gy2 p2 0 y2 0 -0.02
Vsp3 po3 p3 0
Vsr3 p3 pr3 0
Rp3 pr3 0 50
Ru3 u3 0 50
Fr3 u3 0 Vsr3 -1
Fu3 u3 0 Vsp3 -1
Ry3 y3 0 1
Gy3 p3 0 y3 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 4.71114172735079
Cx1 x1 xm1 4.30686999129145e-12
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.649352987731244
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -3.57114254592561
Cx2 x2 xm2 4.30686999129145e-12
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 2.31893208181095
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 0.603618248236217
Cx3 x3 xm3 8.05342537957096e-12
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -0.315251175297791
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -14.2508781347496
Cx4 x4 xm4 8.05342537957096e-12
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 4.49260608100539
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 67.5629168242984
Cx5 x5 xm5 2.88356300968449e-14
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -6.73088179146205e-09
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -9473.92533813877
Cx6 x6 xm6 2.88356300968449e-14
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 6.37678715521492e-05
Rx7 x7 0 1
Fxc7_8 x7 0 Vx8 22755.1998063158
Cx7 x7 xm7 3.27807622205493e-15
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 -9.07782014041513e-10
Rx8 x8 0 1
Fxc8_7 x8 0 Vx7 -2258.54379708303
Cx8 x8 xm8 3.27807622205493e-15
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 2.050265436917e-06
Rx9 x9 0 1
Fxc9_10 x9 0 Vx10 315.517249903735
Cx9 x9 xm9 8.61037113698984e-14
Vx9 xm9 0 0
Gx9_1 x9 0 u1 0 -4.82889560346781e-07
Rx10 x10 0 1
Fxc10_9 x10 0 Vx9 -241.372240484605
Cx10 x10 xm10 8.61037113698984e-14
Vx10 xm10 0 0
Gx10_1 x10 0 u1 0 0.000116556135087528
Rx11 x11 0 1
Fxc11_12 x11 0 Vx12 3473.74789179793
Cx11 x11 xm11 7.36385701297364e-14
Vx11 xm11 0 0
Gx11_1 x11 0 u1 0 -4.30351942173622e-07
Rx12 x12 0 1
Fxc12_11 x12 0 Vx11 -30.4815155248068
Cx12 x12 xm12 7.36385701297364e-14
Vx12 xm12 0 0
Gx12_1 x12 0 u1 0 1.3117779406496e-05
Rx13 x13 0 1
Fxc13_14 x13 0 Vx14 327.588383248525
Cx13 x13 xm13 2.83512527353486e-14
Vx13 xm13 0 0
Gx13_1 x13 0 u1 0 -1.42533797684621e-08
Rx14 x14 0 1
Fxc14_13 x14 0 Vx13 -2258.32542799717
Cx14 x14 xm14 2.83512527353486e-14
Vx14 xm14 0 0
Gx14_1 x14 0 u1 0 3.21887699660183e-05
Rx15 x15 0 1
Fxc15_16 x15 0 Vx16 5.9768606819774
Cx15 x15 xm15 2.47015112633796e-12
Vx15 xm15 0 0
Gx15_1 x15 0 u1 0 -0.00377920994631216
Rx16 x16 0 1
Fxc16_15 x16 0 Vx15 -18.8534512547498
Cx16 x16 xm16 2.47015112633796e-12
Vx16 xm16 0 0
Gx16_1 x16 0 u1 0 0.071251150504262
Rx17 x17 0 1
Fxc17_18 x17 0 Vx18 444.608688899593
Cx17 x17 xm17 6.21082676967847e-14
Vx17 xm17 0 0
Gx17_1 x17 0 u1 0 -1.46135368483712e-07
Rx18 x18 0 1
Fxc18_17 x18 0 Vx17 -359.77972226872
Cx18 x18 xm18 6.21082676967847e-14
Vx18 xm18 0 0
Gx18_1 x18 0 u1 0 5.25765422867068e-05
Rx19 x19 0 1
Fxc19_20 x19 0 Vx20 993.909133806365
Cx19 x19 xm19 6.88618151548846e-14
Vx19 xm19 0 0
Gx19_1 x19 0 u1 0 -2.14454662357434e-07
Rx20 x20 0 1
Fxc20_19 x20 0 Vx19 -135.937236382723
Cx20 x20 xm20 6.88618151548846e-14
Vx20 xm20 0 0
Gx20_1 x20 0 u1 0 2.91523741302595e-05
Rx21 x21 0 1
Fxc21_22 x21 0 Vx22 4276.53551203196
Cx21 x21 xm21 5.46774161318971e-15
Vx21 xm21 0 0
Gx21_1 x21 0 u1 0 -1.47281605630557e-09
Rx22 x22 0 1
Fxc22_21 x22 0 Vx21 -5117.66395969694
Cx22 x22 xm22 5.46774161318971e-15
Vx22 xm22 0 0
Gx22_1 x22 0 u1 0 7.53737765061797e-06
Rx23 x23 0 1
Fxc23_24 x23 0 Vx24 74.6693111994835
Cx23 x23 xm23 1.19014549350492e-13
Vx23 xm23 0 0
Gx23_1 x23 0 u1 0 -2.6261062088855e-07
Rx24 x24 0 1
Fxc24_23 x24 0 Vx23 -634.363023123572
Cx24 x24 xm24 1.19014549350492e-13
Vx24 xm24 0 0
Gx24_1 x24 0 u1 0 0.000166590467371219
Rx25 x25 0 1
Fxc25_26 x25 0 Vx26 25.9333848158752
Cx25 x25 xm25 3.39580797038266e-13
Vx25 xm25 0 0
Gx25_1 x25 0 u1 0 -5.11522220195801e-06
Rx26 x26 0 1
Fxc26_25 x26 0 Vx25 -233.161554780615
Cx26 x26 xm26 3.39580797038266e-13
Vx26 xm26 0 0
Gx26_1 x26 0 u1 0 0.00119267316165685
Rx27 x27 0 1
Fxc27_28 x27 0 Vx28 1425.56447902026
Cx27 x27 xm27 1.0660761974355e-13
Vx27 xm27 0 0
Gx27_1 x27 0 u1 0 -6.51074112680583e-07
Rx28 x28 0 1
Fxc28_27 x28 0 Vx27 -43.5483643821817
Cx28 x28 xm28 1.0660761974355e-13
Vx28 xm28 0 0
Gx28_1 x28 0 u1 0 2.83532126988196e-05
Rx29 x29 0 1
Fxc29_30 x29 0 Vx30 1214.65016289427
Cx29 x29 xm29 6.29358278007233e-14
Vx29 xm29 0 0
Gx29_1 x29 0 u1 0 -1.15888576439023e-07
Rx30 x30 0 1
Fxc30_29 x30 0 Vx29 -153.769733129738
Cx30 x30 xm30 6.29358278007233e-14
Vx30 xm30 0 0
Gx30_1 x30 0 u1 0 1.78201554718137e-05
Rx31 x31 0 1
Fxc31_32 x31 0 Vx32 98.3547331226706
Cx31 x31 xm31 6.18092938643569e-14
Vx31 xm31 0 0
Gx31_1 x31 0 u1 0 -2.73757073847904e-08
Rx32 x32 0 1
Fxc32_31 x32 0 Vx31 -2055.79491547441
Cx32 x32 xm32 6.18092938643569e-14
Vx32 xm32 0 0
Gx32_1 x32 0 u1 0 5.62788400491673e-05
Rx33 x33 0 1
Fxc33_34 x33 0 Vx34 1675.35839816235
Cx33 x33 xm33 5.92714932806977e-14
Vx33 xm33 0 0
Gx33_1 x33 0 u1 0 -1.13622330407649e-07
Rx34 x34 0 1
Fxc34_33 x34 0 Vx33 -137.031095613401
Cx34 x34 xm34 5.92714932806977e-14
Vx34 xm34 0 0
Gx34_1 x34 0 u1 0 1.5569792421908e-05
Rx35 x35 0 1
Fxc35_36 x35 0 Vx36 33.0151596746313
Cx35 x35 xm35 4.85449289847599e-13
Vx35 xm35 0 0
Gx35_1 x35 0 u1 0 -1.17047436733959e-05
Rx36 x36 0 1
Fxc36_35 x36 0 Vx35 -106.337801837521
Cx36 x36 xm36 4.85449289847599e-13
Vx36 xm36 0 0
Gx36_1 x36 0 u1 0 0.00124465671330055
Rx37 x37 0 1
Fxc37_38 x37 0 Vx38 69.4562536856763
Cx37 x37 xm37 7.07373676456137e-14
Vx37 xm37 0 0
Gx37_1 x37 0 u1 0 -2.93634928477335e-08
Rx38 x38 0 1
Fxc38_37 x38 0 Vx37 -2374.10577807345
Cx38 x38 xm38 7.07373676456137e-14
Vx38 xm38 0 0
Gx38_1 x38 0 u1 0 6.97120380342226e-05
Rx39 x39 0 1
Fxc39_40 x39 0 Vx40 155.974759468003
Cx39 x39 xm39 4.92699889036898e-14
Vx39 xm39 0 0
Gx39_1 x39 0 u1 0 -1.67256827843119e-08
Rx40 x40 0 1
Fxc40_39 x40 0 Vx39 -2283.38458348663
Cx40 x40 xm40 4.92699889036898e-14
Vx40 xm40 0 0
Gx40_1 x40 0 u1 0 3.81911662179854e-05
Rx41 x41 0 1
Fxc41_42 x41 0 Vx42 1066.65282285635
Cx41 x41 xm41 1.55367016383078e-13
Vx41 xm41 0 0
Gx41_1 x41 0 u1 0 -5.78013008141146e-07
Rx42 x42 0 1
Fxc42_41 x42 0 Vx41 -34.7391223082737
Cx42 x42 xm42 1.55367016383078e-13
Vx42 xm42 0 0
Gx42_1 x42 0 u1 0 2.00796645855884e-05
Rx43 x43 0 1
Fxc43_44 x43 0 Vx44 69.4666860648144
Cx43 x43 xm43 8.2745464547176e-14
Vx43 xm43 0 0
Gx43_1 x43 0 u1 0 -2.85194132454095e-08
Rx44 x44 0 1
Fxc44_43 x44 0 Vx43 -1960.84772036475
Cx44 x44 xm44 8.2745464547176e-14
Vx44 xm44 0 0
Gx44_1 x44 0 u1 0 5.59222264484014e-05
Rx45 x45 0 1
Fxc45_46 x45 0 Vx46 12.6807677856508
Cx45 x45 xm45 1.78520263333676e-13
Vx45 xm45 0 0
Gx45_1 x45 0 u1 0 -9.19159698150352e-08
Rx46 x46 0 1
Fxc46_45 x46 0 Vx45 -2377.51358939125
Cx46 x46 xm46 1.78520263333676e-13
Vx46 xm46 0 0
Gx46_1 x46 0 u1 0 0.000218531467317322
Rx47 x47 0 1
Fxc47_48 x47 0 Vx48 536.436806250019
Cx47 x47 xm47 1.06144284233908e-13
Vx47 xm47 0 0
Gx47_1 x47 0 u1 0 -2.27376774049975e-07
Rx48 x48 0 1
Fxc48_47 x48 0 Vx47 -161.67839283025
Cx48 x48 xm48 1.06144284233908e-13
Vx48 xm48 0 0
Gx48_1 x48 0 u1 0 3.67619113953269e-05
Rx49 x49 0 1
Fxc49_50 x49 0 Vx50 0.356377512357627
Cx49 x49 xm49 4.03773986408564e-11
Vx49 xm49 0 0
Gx49_1 x49 0 u1 0 -28.8539457384735
Rx50 x50 0 1
Fxc50_49 x50 0 Vx49 -0.563185351774341
Cx50 x50 xm50 4.03773986408564e-11
Vx50 xm50 0 0
Gx50_1 x50 0 u1 0 16.2501195807999
Rx51 x51 0 1
Fxc51_52 x51 0 Vx52 536.461912694153
Cx51 x51 xm51 4.28734109622567e-14
Vx51 xm51 0 0
Gx51_1 x51 0 u1 0 -2.24773653895234e-08
Rx52 x52 0 1
Fxc52_51 x52 0 Vx51 -1026.98008606772
Cx52 x52 xm52 4.28734109622567e-14
Vx52 xm52 0 0
Gx52_1 x52 0 u1 0 2.30838066423082e-05
Rx53 x53 0 1
Fxc53_54 x53 0 Vx54 1047.89565471436
Cx53 x53 xm53 3.84734228551787e-14
Vx53 xm53 0 0
Gx53_1 x53 0 u1 0 -1.85888872893405e-08
Rx54 x54 0 1
Fxc54_53 x54 0 Vx53 -681.474901462236
Cx54 x54 xm54 3.84734228551787e-14
Vx54 xm54 0 0
Gx54_1 x54 0 u1 0 1.2667860133796e-05
Rx55 x55 0 1
Fxc55_56 x55 0 Vx56 12.0826142087576
Cx55 x55 xm55 2.41483364210631e-12
Vx55 xm55 0 0
Gx55_1 x55 0 u1 0 -0.00100242657751205
Rx56 x56 0 1
Fxc56_55 x56 0 Vx55 -15.9638530935828
Cx56 x56 xm56 2.41483364210631e-12
Vx56 xm56 0 0
Gx56_1 x56 0 u1 0 0.0160025906205054
Rx57 x57 0 1
Fxc57_58 x57 0 Vx58 15.535530622417
Cx57 x57 xm57 3.4976618046498e-13
Vx57 xm57 0 0
Gx57_1 x57 0 u1 0 -5.18551892121921e-07
Rx58 x58 0 1
Fxc58_57 x58 0 Vx57 -578.273951913939
Cx58 x58 xm58 3.4976618046498e-13
Vx58 xm58 0 0
Gx58_1 x58 0 u1 0 0.000299865051929794
Rx59 x59 0 1
Fxc59_60 x59 0 Vx60 591.420627989866
Cx59 x59 xm59 1.82634891235488e-14
Vx59 xm59 0 0
Gx59_1 x59 0 u1 0 -1.12494871636132e-09
Rx60 x60 0 1
Fxc60_59 x60 0 Vx59 -5706.09619031033
Cx60 x60 xm60 1.82634891235488e-14
Vx60 xm60 0 0
Gx60_1 x60 0 u1 0 6.41906558472383e-06
Rx61 x61 0 1
Fxc61_62 x61 0 Vx62 1274.12255936988
Cx61 x61 xm61 8.73129447755975e-14
Vx61 xm61 0 0
Gx61_1 x61 0 u1 0 -8.68114207074114e-08
Rx62 x62 0 1
Fxc62_61 x62 0 Vx61 -120.877542143541
Cx62 x62 xm62 8.73129447755975e-14
Vx62 xm62 0 0
Gx62_1 x62 0 u1 0 1.04935511651008e-05
Rx63 x63 0 1
Fxc63_64 x63 0 Vx64 6.22022062773607
Cx63 x63 xm63 1.19432876562705e-11
Vx63 xm63 0 0
Gx63_1 x63 0 u1 0 -0.343913259888117
Rx64 x64 0 1
Fxc64_63 x64 0 Vx63 -1.75579368499634
Cx64 x64 xm64 1.19432876562705e-11
Vx64 xm64 0 0
Gx64_1 x64 0 u1 0 0.603840729898063
Rx65 x65 0 1
Fxc65_66 x65 0 Vx66 39.6687367560648
Cx65 x65 xm65 2.49726015690021e-13
Vx65 xm65 0 0
Gx65_1 x65 0 u1 0 -3.1648832956867e-07
Rx66 x66 0 1
Fxc66_65 x66 0 Vx65 -495.438702795361
Cx66 x66 xm66 2.49726015690021e-13
Vx66 xm66 0 0
Gx66_1 x66 0 u1 0 0.000156800567451373
Rx67 x67 0 1
Fxc67_68 x67 0 Vx68 1187.5088343608
Cx67 x67 xm67 2.53897718170844e-14
Vx67 xm67 0 0
Gx67_1 x67 0 u1 0 -5.93735470051078e-09
Rx68 x68 0 1
Fxc68_67 x68 0 Vx67 -1635.18684782533
Cx68 x68 xm68 2.53897718170844e-14
Vx68 xm68 0 0
Gx68_1 x68 0 u1 0 9.70868431714915e-06
Rx69 x69 0 1
Fxc69_70 x69 0 Vx70 1.24711865767171
Cx69 x69 xm69 2.12240440031949e-11
Vx69 xm69 0 0
Gx69_1 x69 0 u1 0 -1.79724586738083
Rx70 x70 0 1
Fxc70_69 x70 0 Vx69 -2.86690954620997
Cx70 x70 xm70 2.12240440031949e-11
Vx70 xm70 0 0
Gx70_1 x70 0 u1 0 5.15254133408052
Rx71 x71 0 1
Fxc71_72 x71 0 Vx72 1232.80977536121
Cx71 x71 xm71 1.58125194797678e-13
Vx71 xm71 0 0
Gx71_1 x71 0 u1 0 -3.30548000972376e-07
Rx72 x72 0 1
Fxc72_71 x72 0 Vx71 -42.310403406277
Cx72 x72 xm72 1.58125194797678e-13
Vx72 xm72 0 0
Gx72_1 x72 0 u1 0 1.39856192662797e-05
Rx73 x73 0 1
Fxc73_74 x73 0 Vx74 260.425636576108
Cx73 x73 xm73 2.51123986719261e-13
Vx73 xm73 0 0
Gx73_1 x73 0 u1 0 -1.14632119415174e-06
Rx74 x74 0 1
Fxc74_73 x74 0 Vx73 -83.0062268845765
Cx74 x74 xm74 2.51123986719261e-13
Vx74 xm74 0 0
Gx74_1 x74 0 u1 0 9.51517971243576e-05
Rx75 x75 0 1
Fxc75_76 x75 0 Vx76 1170.00761001182
Cx75 x75 xm75 5.50290062427746e-14
Vx75 xm75 0 0
Gx75_1 x75 0 u1 0 -2.65059024886127e-08
Rx76 x76 0 1
Fxc76_75 x76 0 Vx75 -395.037632798858
Cx76 x76 xm76 5.50290062427746e-14
Vx76 xm76 0 0
Gx76_1 x76 0 u1 0 1.04708289742989e-05
Rx77 x77 0 1
Fxc77_78 x77 0 Vx78 347.701210991986
Cx77 x77 xm77 1.73036537262631e-13
Vx77 xm77 0 0
Gx77_1 x77 0 u1 0 -4.53510705761923e-07
Rx78 x78 0 1
Fxc78_77 x78 0 Vx77 -139.994659286797
Cx78 x78 xm78 1.73036537262631e-13
Vx78 xm78 0 0
Gx78_1 x78 0 u1 0 6.34890767360553e-05
Rx79 x79 0 1
Fxc79_80 x79 0 Vx80 40.1836295673689
Cx79 x79 xm79 1.04005943428604e-12
Vx79 xm79 0 0
Gx79_1 x79 0 u1 0 -4.55066015076472e-05
Rx80 x80 0 1
Fxc80_79 x80 0 Vx79 -34.3314249452786
Cx80 x80 xm80 1.04005943428604e-12
Vx80 xm80 0 0
Gx80_1 x80 0 u1 0 0.00156230647417449
Rx81 x81 0 1
Fxc81_82 x81 0 Vx82 44.3006273057236
Cx81 x81 xm81 1.69597975933452e-13
Vx81 xm81 0 0
Gx81_1 x81 0 u1 0 -7.50142769424825e-08
Rx82 x82 0 1
Fxc82_81 x82 0 Vx81 -1197.04118441021
Cx82 x82 xm82 1.69597975933451e-13
Vx82 xm82 0 0
Gx82_1 x82 0 u1 0 8.97951789189048e-05
Rx83 x83 0 1
Fxc83_84 x83 0 Vx84 1341.34590783269
Cx83 x83 xm83 1.6574520023931e-13
Vx83 xm83 0 0
Gx83_1 x83 0 u1 0 -3.3176229131289e-07
Rx84 x84 0 1
Fxc84_83 x84 0 Vx83 -43.2176385575793
Cx84 x84 xm84 1.6574520023931e-13
Vx84 xm84 0 0
Gx84_1 x84 0 u1 0 1.43379827929948e-05
Rx85 x85 0 1
Fxc85_86 x85 0 Vx86 121.87279599379
Cx85 x85 xm85 4.17930149743441e-14
Vx85 xm85 0 0
Gx85_1 x85 0 u1 0 -1.47312415497432e-09
Rx86 x86 0 1
Fxc86_85 x86 0 Vx85 -7847.20405058023
Cx86 x86 xm86 4.17930149743441e-14
Vx86 xm86 0 0
Gx86_1 x86 0 u1 0 1.15599058359221e-05
Rx87 x87 0 1
Fxc87_88 x87 0 Vx88 353.375902372115
Cx87 x87 xm87 9.47540753730688e-14
Vx87 xm87 0 0
Gx87_1 x87 0 u1 0 -5.03336697572282e-08
Rx88 x88 0 1
Fxc88_87 x88 0 Vx87 -542.31590753162
Cx88 x88 xm88 9.47540753730688e-14
Vx88 xm88 0 0
Gx88_1 x88 0 u1 0 2.72967497937881e-05
Rx89 x89 0 1
Fxc89_90 x89 0 Vx90 134.687710616814
Cx89 x89 xm89 3.39327012867075e-13
Vx89 xm89 0 0
Gx89_1 x89 0 u1 0 -8.69256001869561e-07
Rx90 x90 0 1
Fxc90_89 x90 0 Vx89 -114.855215852665
Cx90 x90 xm90 3.39327012867075e-13
Vx90 xm90 0 0
Gx90_1 x90 0 u1 0 9.98385857259532e-05
Rx91 x91 0 1
Fxc91_92 x91 0 Vx92 1394.96654096327
Cx91 x91 xm91 2.21690564685036e-14
Vx91 xm91 0 0
Gx91_1 x91 0 u1 0 -3.97442485099303e-09
Rx92 x92 0 1
Fxc92_91 x92 0 Vx91 -2671.26647259847
Cx92 x92 xm92 2.21690564685036e-14
Vx92 xm92 0 0
Gx92_1 x92 0 u1 0 1.06167478523199e-05
Rx93 x93 0 1
Fxc93_94 x93 0 Vx94 1146.52430229269
Cx93 x93 xm93 1.4311943973241e-13
Vx93 xm93 0 0
Gx93_1 x93 0 u1 0 -1.18741515724191e-07
Rx94 x94 0 1
Fxc94_93 x94 0 Vx93 -82.2503523738923
Cx94 x94 xm94 1.4311943973241e-13
Vx94 xm94 0 0
Gx94_1 x94 0 u1 0 9.76653150972482e-06
Rx95 x95 0 1
Fxc95_96 x95 0 Vx96 152.52342999519
Cx95 x95 xm95 1.49527034425067e-14
Vx95 xm95 0 0
Gx95_1 x95 0 u1 0 -2.75125506761358e-10
Rx96 x96 0 1
Fxc96_95 x96 0 Vx95 -59050.4255701591
Cx96 x96 xm96 1.49527034425067e-14
Vx96 xm96 0 0
Gx96_1 x96 0 u1 0 1.62462782594639e-05
Rx97 x97 0 1
Fxc97_98 x97 0 Vx98 65.1316295382976
Cx97 x97 xm97 1.29249231176747e-13
Vx97 xm97 0 0
Gx97_1 x97 0 u1 0 -1.8773255377285e-08
Rx98 x98 0 1
Fxc98_97 x98 0 Vx97 -1921.27591327259
Cx98 x98 xm98 1.29249231176747e-13
Vx98 xm98 0 0
Gx98_1 x98 0 u1 0 3.6068603370093e-05
Rx99 x99 0 1
Fxc99_100 x99 0 Vx100 1523.11400961381
Cx99 x99 xm99 2.97577142965506e-14
Vx99 xm99 0 0
Gx99_1 x99 0 u1 0 -6.7805459020016e-09
Rx100 x100 0 1
Fxc100_99 x100 0 Vx99 -1608.84998836577
Cx100 x100 xm100 2.97577142965506e-14
Vx100 xm100 0 0
Gx100_1 x100 0 u1 0 1.09088811955488e-05
Rx101 x101 0 1
Fxc101_102 x101 0 Vx102 173.454675830585
Cx101 x101 xm101 3.66480875628994e-13
Vx101 xm101 0 0
Gx101_1 x101 0 u1 0 -6.51466093981107e-07
Rx102 x102 0 1
Fxc102_101 x102 0 Vx101 -96.544306679683
Cx102 x102 xm102 3.66480875628994e-13
Vx102 xm102 0 0
Gx102_1 x102 0 u1 0 6.28953423687272e-05
Rx103 x103 0 1
Fxc103_104 x103 0 Vx104 1109.24735846092
Cx103 x103 xm103 1.55725403798337e-13
Vx103 xm103 0 0
Gx103_1 x103 0 u1 0 -1.24153138361159e-07
Rx104 x104 0 1
Fxc104_103 x104 0 Vx103 -87.1394331375762
Cx104 x104 xm104 1.55725403798337e-13
Vx104 xm104 0 0
Gx104_1 x104 0 u1 0 1.08186340990425e-05
Rx105 x105 0 1
Fxc105_106 x105 0 Vx106 1472.9406610034
Cx105 x105 xm105 2.70690945024366e-14
Vx105 xm105 0 0
Gx105_1 x105 0 u1 0 -4.07705863309248e-09
Rx106 x106 0 1
Fxc106_105 x106 0 Vx105 -2383.14014593404
Cx106 x106 xm106 2.70690945024366e-14
Vx106 xm106 0 0
Gx106_1 x106 0 u1 0 9.71620210584966e-06
Rx107 x107 0 1
Fxc107_108 x107 0 Vx108 4189.51073694025
Cx107 x107 xm107 1.05947857159888e-13
Vx107 xm107 0 0
Gx107_1 x107 0 u1 0 -6.55689986649896e-08
Rx108 x108 0 1
Fxc108_107 x108 0 Vx107 -52.483624398605
Cx108 x108 xm108 1.05947857159888e-13
Vx108 xm108 0 0
Gx108_1 x108 0 u1 0 3.44129869812595e-06
Rx109 x109 0 1
Fxc109_110 x109 0 Vx110 1449.48530620349
Cx109 x109 xm109 8.05411899100067e-14
Vx109 xm109 0 0
Gx109_1 x109 0 u1 0 -3.47738716289156e-08
Rx110 x110 0 1
Fxc110_109 x110 0 Vx109 -292.580822253074
Cx110 x110 xm110 8.05411899100067e-14
Vx110 xm110 0 0
Gx110_1 x110 0 u1 0 1.0174167954111e-05
Rx111 x111 0 1
Fxc111_112 x111 0 Vx112 350.194109912843
Cx111 x111 xm111 2.77463484357731e-13
Vx111 xm111 0 0
Gx111_1 x111 0 u1 0 -2.59376256859559e-07
Rx112 x112 0 1
Fxc112_111 x112 0 Vx111 -105.682742565954
Cx112 x112 xm112 2.77463484357731e-13
Vx112 xm112 0 0
Gx112_1 x112 0 u1 0 2.74115941814094e-05
Rx113 x113 0 1
Cx113 x113 0 1.26327330229509e-10
Gx113_1 x113 0 u1 0 -5.2482619018823
Rx114 x114 0 1
Fxc114_115 x114 0 Vx115 1179.66817957751
Cx114 x114 xm114 1.99280702854811e-13
Vx114 xm114 0 0
Gx114_1 x114 0 u1 0 -2.51065931436558e-07
Rx115 x115 0 1
Fxc115_114 x115 0 Vx114 -63.6651141382228
Cx115 x115 xm115 1.99280702854811e-13
Vx115 xm115 0 0
Gx115_1 x115 0 u1 0 1.59841411811277e-05
Rx116 x116 0 1
Fxc116_117 x116 0 Vx117 816.072477240114
Cx116 x116 xm116 3.34725367390173e-14
Vx116 xm116 0 0
Gx116_1 x116 0 u1 0 -3.36089290178885e-09
Rx117 x117 0 1
Fxc117_116 x117 0 Vx116 -3443.35930131658
Cx117 x117 xm117 3.34725367390174e-14
Vx117 xm117 0 0
Gx117_1 x117 0 u1 0 1.15727618341035e-05
Rx118 x118 0 1
Fxc118_119 x118 0 Vx119 66.2203039474744
Cx118 x118 xm118 1.20981905835219e-12
Vx118 xm118 0 0
Gx118_1 x118 0 u1 0 -1.18221794985669e-05
Rx119 x119 0 1
Fxc119_118 x119 0 Vx118 -33.5655137123057
Cx119 x119 xm119 1.20981905835219e-12
Vx119 xm119 0 0
Gx119_1 x119 0 u1 0 0.000396817528068487
Rx120 x120 0 1
Fxc120_121 x120 0 Vx121 32.8189478591376
Cx120 x120 xm120 2.41747187333388e-13
Vx120 xm120 0 0
Gx120_1 x120 0 u1 0 -4.78840791907876e-08
Rx121 x121 0 1
Fxc121_120 x121 0 Vx120 -1833.79003669021
Cx121 x121 xm121 2.41747187333388e-13
Vx121 xm121 0 0
Gx121_1 x121 0 u1 0 8.78093473361514e-05
Rx122 x122 0 1
Fxc122_123 x122 0 Vx123 87.0483224959785
Cx122 x122 xm122 6.05595987313277e-13
Vx122 xm122 0 0
Gx122_1 x122 0 u1 0 -1.76604882800903e-06
Rx123 x123 0 1
Fxc123_122 x123 0 Vx122 -112.677776245508
Cx123 x123 xm123 6.05595987313277e-13
Vx123 xm123 0 0
Gx123_1 x123 0 u1 0 0.000198994454681044
Rx124 x124 0 1
Fxc124_125 x124 0 Vx125 8.34985941078969
Cx124 x124 xm124 4.27273098109608e-12
Vx124 xm124 0 0
Gx124_1 x124 0 u1 0 -0.000361725499489477
Rx125 x125 0 1
Fxc125_124 x125 0 Vx124 -27.5794889153617
Cx125 x125 xm125 4.27273098109608e-12
Vx125 xm125 0 0
Gx125_1 x125 0 u1 0 0.0099762044035737
Rx126 x126 0 1
Fxc126_127 x126 0 Vx127 1373.73381840876
Cx126 x126 xm126 2.2113064440014e-13
Vx126 xm126 0 0
Gx126_1 x126 0 u1 0 -2.45853519237459e-07
Rx127 x127 0 1
Fxc127_126 x127 0 Vx126 -58.1632040134788
Cx127 x127 xm127 2.2113064440014e-13
Vx127 xm127 0 0
Gx127_1 x127 0 u1 0 1.42996283968401e-05
Rx128 x128 0 1
Fxc128_129 x128 0 Vx129 19.3461561044746
Cx128 x128 xm128 3.84635353963742e-13
Vx128 xm128 0 0
Gx128_1 x128 0 u1 0 -9.28328055530745e-08
Rx129 x129 0 1
Fxc129_128 x129 0 Vx128 -1434.03122010332
Cx129 x129 xm129 3.84635353963742e-13
Vx129 xm129 0 0
Gx129_1 x129 0 u1 0 0.00013312514141289
Rx130 x130 0 1
Fxc130_131 x130 0 Vx131 10.7270261935519
Cx130 x130 xm130 1.31174697600352e-12
Vx130 xm130 0 0
Gx130_1 x130 0 u1 0 -8.3035638841843e-06
Rx131 x131 0 1
Fxc131_130 x131 0 Vx130 -236.31045724118
Cx131 x131 xm131 1.31174697600352e-12
Vx131 xm131 0 0
Gx131_1 x131 0 u1 0 0.00196221897820294
Rx132 x132 0 1
Fxc132_133 x132 0 Vx133 377.402009568768
Cx132 x132 xm132 6.73245820833979e-13
Vx132 xm132 0 0
Gx132_1 x132 0 u1 0 -4.48036811381799e-06
Rx133 x133 0 1
Fxc133_132 x133 0 Vx132 -25.9472222942777
Cx133 x133 xm133 6.73245820833979e-13
Vx133 xm133 0 0
Gx133_1 x133 0 u1 0 0.000116253107409429
Rx134 x134 0 1
Fxc134_135 x134 0 Vx135 232.758352553756
Cx134 x134 xm134 5.84808784752663e-13
Vx134 xm134 0 0
Gx134_1 x134 0 u1 0 -1.29389080399073e-06
Rx135 x135 0 1
Fxc135_134 x135 0 Vx134 -61.4626990398924
Cx135 x135 xm135 5.84808784752663e-13
Vx135 xm135 0 0
Gx135_1 x135 0 u1 0 7.95260210761665e-05
Rx136 x136 0 1
Fxc136_137 x136 0 Vx137 207.141788705059
Cx136 x136 xm136 1.79416446898388e-13
Vx136 xm136 0 0
Gx136_1 x136 0 u1 0 -2.18726982435231e-08
Rx137 x137 0 1
Fxc137_136 x137 0 Vx136 -801.435551699879
Cx137 x137 xm137 1.79416446898388e-13
Vx137 xm137 0 0
Gx137_1 x137 0 u1 0 1.75295579839629e-05
Rx138 x138 0 1
Fxc138_139 x138 0 Vx139 181.127379569173
Cx138 x138 xm138 9.55321996041439e-13
Vx138 xm138 0 0
Gx138_1 x138 0 u1 0 -3.37061150756012e-06
Rx139 x139 0 1
Fxc139_138 x139 0 Vx138 -35.3223174847751
Cx139 x139 xm139 9.55321996041439e-13
Vx139 xm139 0 0
Gx139_1 x139 0 u1 0 0.000119057809787875
Rx140 x140 0 1
Fxc140_141 x140 0 Vx141 23.1933332113227
Cx140 x140 xm140 4.22656817502044e-13
Vx140 xm140 0 0
Gx140_1 x140 0 u1 0 -6.15450144654684e-08
Rx141 x141 0 1
Fxc141_140 x141 0 Vx140 -1459.66127742099
Cx141 x141 xm141 4.22656817502044e-13
Vx141 xm141 0 0
Gx141_1 x141 0 u1 0 8.98348744335592e-05
Rx142 x142 0 1
Fxc142_143 x142 0 Vx143 61.2300859783102
Cx142 x142 xm142 2.32688864615857e-12
Vx142 xm142 0 0
Gx142_1 x142 0 u1 0 -2.29189079276921e-05
Rx143 x143 0 1
Fxc143_142 x143 0 Vx142 -20.005110738955
Cx143 x143 xm143 2.32688864615857e-12
Vx143 xm143 0 0
Gx143_1 x143 0 u1 0 0.000458495291109394
Rx144 x144 0 1
Fxc144_145 x144 0 Vx145 557.560547924165
Cx144 x144 xm144 2.24826805546157e-13
Vx144 xm144 0 0
Gx144_1 x144 0 u1 0 -9.94221123212158e-08
Rx145 x145 0 1
Fxc145_144 x145 0 Vx144 -236.36060215471
Cx145 x145 xm145 2.24826805546157e-13
Vx145 xm145 0 0
Gx145_1 x145 0 u1 0 2.34994703357358e-05
Rx146 x146 0 1
Fxc146_147 x146 0 Vx147 436.944480191724
Cx146 x146 xm146 7.62490228495289e-13
Vx146 xm146 0 0
Gx146_1 x146 0 u1 0 -9.40774372228672e-07
Rx147 x147 0 1
Fxc147_146 x147 0 Vx146 -29.6840505017269
Cx147 x147 xm147 7.62490228495289e-13
Vx147 xm147 0 0
Gx147_1 x147 0 u1 0 2.79259939759663e-05
Rx148 x148 0 1
Fxc148_149 x148 0 Vx149 42.0746481549003
Cx148 x148 xm148 3.12815339647046e-13
Vx148 xm148 0 0
Gx148_1 x148 0 u1 0 -2.41001633908674e-08
Rx149 x149 0 1
Fxc149_148 x149 0 Vx148 -1993.63724371182
Cx149 x149 xm149 3.12815339647046e-13
Vx149 xm149 0 0
Gx149_1 x149 0 u1 0 4.80469833155735e-05
Rx150 x150 0 1
Fxc150_151 x150 0 Vx151 11.2679580764121
Cx150 x150 xm150 1.21980473796757e-12
Vx150 xm150 0 0
Gx150_1 x150 0 u1 0 -4.40817784454114e-07
Rx151 x151 0 1
Fxc151_150 x151 0 Vx150 -514.060668532967
Cx151 x151 xm151 1.21980473796757e-12
Vx151 xm151 0 0
Gx151_1 x151 0 u1 0 0.000226607084977703
Rx152 x152 0 1
Fxc152_153 x152 0 Vx153 2.80486045794338
Cx152 x152 xm152 6.30927595670662e-12
Vx152 xm152 0 0
Gx152_1 x152 0 u1 0 -4.60035744654429e-05
Rx153 x153 0 1
Fxc153_152 x153 0 Vx152 -91.255538481971
Cx153 x153 xm153 6.30927595670662e-12
Vx153 xm153 0 0
Gx153_1 x153 0 u1 0 0.00419808095993944
Rx154 x154 0 1
Fxc154_155 x154 0 Vx155 7419.62081704781
Cx154 x154 xm154 5.94898906330198e-14
Vx154 xm154 0 0
Gx154_1 x154 0 u1 0 -1.1663864474428e-08
Rx155 x155 0 1
Fxc155_154 x155 0 Vx154 -379.892945902257
Cx155 x155 xm155 5.94898906330198e-14
Vx155 xm155 0 0
Gx155_1 x155 0 u1 0 4.43101983579512e-06
Rx156 x156 0 1
Fxc156_157 x156 0 Vx157 609.587040127488
Cx156 x156 xm156 1.88629779420802e-12
Vx156 xm156 0 0
Gx156_1 x156 0 u1 0 -9.98305095575484e-06
Rx157 x157 0 1
Fxc157_156 x157 0 Vx156 -5.03287207985895
Cx157 x157 xm157 1.88629779420802e-12
Vx157 xm157 0 0
Gx157_1 x157 0 u1 0 5.02434184270277e-05
Rx158 x158 0 1
Fxc158_159 x158 0 Vx159 15.7096826799385
Cx158 x158 xm158 2.53255697284169e-12
Vx158 xm158 0 0
Gx158_1 x158 0 u1 0 -5.64532129840827e-06
Rx159 x159 0 1
Fxc159_158 x159 0 Vx158 -127.443108417839
Cx159 x159 xm159 2.53255697284169e-12
Vx159 xm159 0 0
Gx159_1 x159 0 u1 0 0.00071945729428658
Rx160 x160 0 1
Fxc160_161 x160 0 Vx161 25.4723146587905
Cx160 x160 xm160 1.07068178225324e-12
Vx160 xm160 0 0
Gx160_1 x160 0 u1 0 -4.28548305936242e-07
Rx161 x161 0 1
Fxc161_160 x161 0 Vx160 -470.125188941025
Cx161 x161 xm161 1.07068178225324e-12
Vx161 xm161 0 0
Gx161_1 x161 0 u1 0 0.000201471353298632
Rx162 x162 0 1
Cx162 x162 0 5.22190407222509e-10
Gx162_1 x162 0 u1 0 -0.866840315988095
Rx163 x163 0 1
Fxc163_164 x163 0 Vx164 180.08518240188
Cx163 x163 xm163 1.10121754249303e-12
Vx163 xm163 0 0
Gx163_1 x163 0 u1 0 -7.59604906106668e-07
Rx164 x164 0 1
Fxc164_163 x164 0 Vx163 -76.5627990474259
Cx164 x164 xm164 1.10121754249303e-12
Vx164 xm164 0 0
Gx164_1 x164 0 u1 0 5.81574777816836e-05
Rx165 x165 0 1
Fxc165_166 x165 0 Vx166 128.418468643151
Cx165 x165 xm165 1.3584005978461e-12
Vx165 xm165 0 0
Gx165_1 x165 0 u1 0 -1.20483527836428e-06
Rx166 x166 0 1
Fxc166_165 x166 0 Vx165 -80.6291573613597
Cx166 x166 xm166 1.35840059784609e-12
Vx166 xm166 0 0
Gx166_1 x166 0 u1 0 9.71448532537515e-05
Rx167 x167 0 1
Fxc167_168 x167 0 Vx168 3.46348798495064
Cx167 x167 xm167 1.37582820475616e-11
Vx167 xm167 0 0
Gx167_1 x167 0 u1 0 -0.000109084679455464
Rx168 x168 0 1
Fxc168_167 x168 0 Vx167 -40.2651360874888
Cx168 x168 xm168 1.37582820475616e-11
Vx168 xm168 0 0
Gx168_1 x168 0 u1 0 0.00439230946333437
Rx169 x169 0 1
Fxc169_170 x169 0 Vx170 8.35516441509579
Cx169 x169 xm169 2.55525080407755e-12
Vx169 xm169 0 0
Gx169_1 x169 0 u1 0 -2.2854787950552e-06
Rx170 x170 0 1
Fxc170_169 x170 0 Vx169 -267.109869558875
Cx170 x170 xm170 2.55525080407755e-12
Vx170 xm170 0 0
Gx170_1 x170 0 u1 0 0.00061047394282677
Rx171 x171 0 1
Fxc171_172 x171 0 Vx172 1.58957806884633
Cx171 x171 xm171 3.52048110577458e-12
Vx171 xm171 0 0
Gx171_1 x171 0 u1 0 -4.24554699672007e-07
Rx172 x172 0 1
Fxc172_171 x172 0 Vx171 -1110.57244483831
Cx172 x172 xm172 3.52048110577458e-12
Vx172 xm172 0 0
Gx172_1 x172 0 u1 0 0.000471498750782334
Rx173 x173 0 1
Fxc173_174 x173 0 Vx174 2.9866217307126
Cx173 x173 xm173 8.01925764208566e-11
Vx173 xm173 0 0
Gx173_1 x173 0 u1 0 -0.0230983635326091
Rx174 x174 0 1
Fxc174_173 x174 0 Vx173 -2.61536943758414
Cx174 x174 xm174 8.01925764208566e-11
Vx174 xm174 0 0
Gx174_1 x174 0 u1 0 0.0604107540413939
Rx175 x175 0 1
Fxc175_176 x175 0 Vx176 10.5222198350012
Cx175 x175 xm175 1.34818539204243e-12
Vx175 xm175 0 0
Gx175_1 x175 0 u1 0 -8.81527763721093e-08
Rx176 x176 0 1
Fxc176_175 x176 0 Vx175 -1434.28620527811
Cx176 x176 xm176 1.34818539204243e-12
Vx176 xm176 0 0
Gx176_1 x176 0 u1 0 0.000126436311107482
Rx177 x177 0 1
Fxc177_178 x177 0 Vx178 1.19239294253459
Cx177 x177 xm177 2.60286578934868e-10
Vx177 xm177 0 0
Gx177_1 x177 0 u1 0 -0.0547979827428292
Rx178 x178 0 1
Fxc178_177 x178 0 Vx177 -2.46862514459476
Cx178 x178 xm178 2.60286578934868e-10
Vx178 xm178 0 0
Gx178_1 x178 0 u1 0 0.135275678072018
Rx179 x179 0 1
Fxc179_180 x179 0 Vx180 9.13901176004122
Cx179 x179 xm179 1.94992797826926e-12
Vx179 xm179 0 0
Gx179_1 x179 0 u1 0 -1.38307987887476e-07
Rx180 x180 0 1
Fxc180_179 x180 0 Vx179 -985.264579907437
Cx180 x180 xm180 1.94992797826926e-12
Vx180 xm180 0 0
Gx180_1 x180 0 u1 0 0.000136269961583797
Rx181 x181 0 1
Fxc181_182 x181 0 Vx182 88.7010423069764
Cx181 x181 xm181 2.33413529363335e-12
Vx181 xm181 0 0
Gx181_1 x181 0 u1 0 -3.92322838231253e-07
Rx182 x182 0 1
Fxc182_181 x182 0 Vx181 -184.057054563326
Cx182 x182 xm182 2.33413529363335e-12
Vx182 xm182 0 0
Gx182_1 x182 0 u1 0 7.22097860427686e-05
Rx183 x183 0 1
Fxc183_184 x183 0 Vx184 14.0152950264803
Cx183 x183 xm183 1.72271737747677e-11
Vx183 xm183 0 0
Gx183_1 x183 0 u1 0 -0.000109013010637594
Rx184 x184 0 1
Fxc184_183 x184 0 Vx183 -14.8670846912857
Cx184 x184 xm184 1.72271737747677e-11
Vx184 xm184 0 0
Gx184_1 x184 0 u1 0 0.00162070566160114
Rx185 x185 0 1
Fxc185_186 x185 0 Vx186 275.60216660546
Cx185 x185 xm185 3.38373728470339e-12
Vx185 xm185 0 0
Gx185_1 x185 0 u1 0 -4.07605995395669e-06
Rx186 x186 0 1
Fxc186_185 x186 0 Vx185 -13.5068548165017
Cx186 x186 xm186 3.38373728470339e-12
Vx186 xm186 0 0
Gx186_1 x186 0 u1 0 5.50547500214494e-05
Rx187 x187 0 1
Fxc187_188 x187 0 Vx188 34.2456055011797
Cx187 x187 xm187 5.83456226648167e-12
Vx187 xm187 0 0
Gx187_1 x187 0 u1 0 -1.36632883056912e-06
Rx188 x188 0 1
Fxc188_187 x188 0 Vx187 -124.677196536631
Cx188 x188 xm188 5.83456226648167e-12
Vx188 xm188 0 0
Gx188_1 x188 0 u1 0 0.000170350048142532
Rx189 x189 0 1
Fxc189_190 x189 0 Vx190 38.8233229767543
Cx189 x189 xm189 3.71913677806581e-11
Vx189 xm189 0 0
Gx189_1 x189 0 u1 0 -0.00239702232028316
Rx190 x190 0 1
Fxc190_189 x190 0 Vx189 -4.87584470757265
Cx190 x190 xm190 3.71913677806581e-11
Vx190 xm190 0 0
Gx190_1 x190 0 u1 0 0.0116875085942862
Rx191 x191 0 1
Fxc191_192 x191 0 Vx192 33.5097289105636
Cx191 x191 xm191 3.43647746350443e-11
Vx191 xm191 0 0
Gx191_1 x191 0 u1 0 -0.00188805468748062
Rx192 x192 0 1
Fxc192_191 x192 0 Vx191 -6.58382475058671
Cx192 x192 xm192 3.43647746350443e-11
Vx192 xm192 0 0
Gx192_1 x192 0 u1 0 0.0124306211818961
Rx193 x193 0 1
Fxc193_194 x193 0 Vx194 1.81130733370953
Cx193 x193 xm193 1.92407202503742e-10
Vx193 xm193 0 0
Gx193_1 x193 0 u1 0 -0.000489783018731503
Rx194 x194 0 1
Fxc194_193 x194 0 Vx193 -13.5353249335575
Cx194 x194 xm194 1.92407202503742e-10
Vx194 xm194 0 0
Gx194_1 x194 0 u1 0 0.00662937230546957
Rx195 x195 0 1
Fxc195_196 x195 0 Vx196 217.665581252764
Cx195 x195 xm195 8.89563374249556e-13
Vx195 xm195 0 0
Gx195_1 x195 0 u1 0 -1.01040650699523e-07
Rx196 x196 0 1
Fxc196_195 x196 0 Vx195 -342.516819611612
Cx196 x196 xm196 8.89563374249556e-13
Vx196 xm196 0 0
Gx196_1 x196 0 u1 0 3.46081223290885e-05
Rx197 x197 0 1
Fxc197_198 x197 0 Vx198 1.58251524871887
Cx197 x197 xm197 1.38719414317867e-09
Vx197 xm197 0 0
Gx197_1 x197 0 u1 0 -0.0819647826272169
Rx198 x198 0 1
Fxc198_197 x198 0 Vx197 -0.368098062785082
Cx198 x198 xm198 1.38719414317867e-09
Vx198 xm198 0 0
Gx198_1 x198 0 u1 0 0.0301710777016789
Rx199 x199 0 1
Cx199 x199 0 4.58826427740312e-07
Gx199_1 x199 0 u1 0 -0.664245904842795
Rx200 x200 0 1
Cx200 x200 0 7.53723517430562e-08
Gx200_1 x200 0 u1 0 -0.151468769908563
Rx201 x201 0 1
Fxc201_202 x201 0 Vx202 2.11245107764624
Cx201 x201 xm201 4.30686999129145e-12
Vx201 xm201 0 0
Gx201_2 x201 0 u2 0 -0.0871763805726945
Rx202 x202 0 1
Fxc202_201 x202 0 Vx201 -7.96428321605149
Cx202 x202 xm202 4.30686999129145e-12
Vx202 xm202 0 0
Gx202_2 x202 0 u2 0 0.694297384631228
Rx203 x203 0 1
Fxc203_204 x203 0 Vx204 1.41615349491078
Cx203 x203 xm203 8.05342537957096e-12
Vx203 xm203 0 0
Gx203_2 x203 0 u2 0 -0.112505761797602
Rx204 x204 0 1
Fxc204_203 x204 0 Vx203 -6.0742639314443
Cx204 x204 xm204 8.05342537957096e-12
Vx204 xm204 0 0
Gx204_2 x204 0 u2 0 0.68338969096684
Rx205 x205 0 1
Fxc205_206 x205 0 Vx206 565.62639185662
Cx205 x205 xm205 2.88356300968449e-14
Vx205 xm205 0 0
Gx205_2 x205 0 u2 0 -1.49279908714582e-08
Rx206 x206 0 1
Fxc206_205 x206 0 Vx205 -1131.64102459798
Cx206 x206 xm206 2.88356300968449e-14
Vx206 xm206 0 0
Gx206_2 x206 0 u2 0 1.68931268849662e-05
Rx207 x207 0 1
Fxc207_208 x207 0 Vx208 3410.76409919652
Cx207 x207 xm207 3.27807622205493e-15
Vx207 xm207 0 0
Gx207_2 x207 0 u2 0 -2.32209721388818e-10
Rx208 x208 0 1
Fxc208_207 x208 0 Vx207 -15068.0650667241
Cx208 x208 xm208 3.27807622205493e-15
Vx208 xm208 0 0
Gx208_2 x208 0 u2 0 3.49895119101258e-06
Rx209 x209 0 1
Fxc209_210 x209 0 Vx210 1170.08163988478
Cx209 x209 xm209 8.61037113698984e-14
Vx209 xm209 0 0
Gx209_2 x209 0 u2 0 -1.71512173222054e-07
Rx210 x210 0 1
Fxc210_209 x210 0 Vx209 -65.0870015602543
Cx210 x210 xm210 8.61037113698983e-14
Vx210 xm210 0 0
Gx210_2 x210 0 u2 0 1.11632130861065e-05
Rx211 x211 0 1
Fxc211_212 x211 0 Vx212 371.444525094883
Cx211 x211 xm211 7.36385701297364e-14
Vx211 xm211 0 0
Gx211_2 x211 0 u2 0 -7.21032677085364e-08
Rx212 x212 0 1
Fxc212_211 x212 0 Vx211 -285.063025941911
Cx212 x212 xm212 7.36385701297364e-14
Vx212 xm212 0 0
Gx212_2 x212 0 u2 0 2.05539756732951e-05
Rx213 x213 0 1
Fxc213_214 x213 0 Vx214 844.133729459617
Cx213 x213 xm213 2.83512527353486e-14
Vx213 xm213 0 0
Gx213_2 x213 0 u2 0 -8.26612986238768e-09
Rx214 x214 0 1
Fxc214_213 x214 0 Vx213 -876.402813900375
Cx214 x214 xm214 2.83512527353486e-14
Vx214 xm214 0 0
Gx214_2 x214 0 u2 0 7.24445947146247e-06
Rx215 x215 0 1
Fxc215_216 x215 0 Vx216 11.5698609699591
Cx215 x215 xm215 2.47015112633796e-12
Vx215 xm215 0 0
Gx215_2 x215 0 u2 0 -0.00238477224240134
Rx216 x216 0 1
Fxc216_215 x216 0 Vx215 -9.73948190187202
Cx216 x216 xm216 2.47015112633796e-12
Vx216 xm216 0 0
Gx216_2 x216 0 u2 0 0.0232264460949546
Rx217 x217 0 1
Fxc217_218 x217 0 Vx218 176.912666906066
Cx217 x217 xm217 6.21082676967847e-14
Vx217 xm217 0 0
Gx217_2 x217 0 u2 0 -2.3952910363556e-08
Rx218 x218 0 1
Fxc218_217 x218 0 Vx217 -904.181670018509
Cx218 x218 xm218 6.21082676967847e-14
Vx218 xm218 0 0
Gx218_2 x218 0 u2 0 2.16577824943237e-05
Rx219 x219 0 1
Fxc219_220 x219 0 Vx220 502.932321898951
Cx219 x219 xm219 6.88618151548846e-14
Vx219 xm219 0 0
Gx219_2 x219 0 u2 0 -5.16259486201728e-08
Rx220 x220 0 1
Fxc220_219 x220 0 Vx219 -268.643026073654
Cx220 x220 xm220 6.88618151548846e-14
Vx220 xm220 0 0
Gx220_2 x220 0 u2 0 1.38689510612462e-05
Rx221 x221 0 1
Fxc221_222 x221 0 Vx222 9041.78763180782
Cx221 x221 xm221 5.46774161318971e-15
Vx221 xm221 0 0
Gx221_2 x221 0 u2 0 -5.75626040171615e-10
Rx222 x222 0 1
Fxc222_221 x222 0 Vx221 -2420.52485122504
Cx222 x222 xm222 5.46774161318971e-15
Vx222 xm222 0 0
Gx222_2 x222 0 u2 0 1.39331713524766e-06
Rx223 x223 0 1
Fxc223_224 x223 0 Vx224 268.519773184137
Cx223 x223 xm223 1.19014549350492e-13
Vx223 xm223 0 0
Gx223_2 x223 0 u2 0 -1.74325577643665e-07
Rx224 x224 0 1
Fxc224_223 x224 0 Vx223 -176.402092945971
Cx224 x224 xm224 1.19014549350492e-13
Vx224 xm224 0 0
Gx224_2 x224 0 u2 0 3.07513967503579e-05
Rx225 x225 0 1
Fxc225_226 x225 0 Vx226 113.164811409368
Cx225 x225 xm225 3.39580797038266e-13
Vx225 xm225 0 0
Gx225_2 x225 0 u2 0 -2.93827354061806e-06
Rx226 x226 0 1
Fxc226_225 x226 0 Vx225 -53.432407557504
Cx226 x226 xm226 3.39580797038266e-13
Vx226 xm226 0 0
Gx226_2 x226 0 u2 0 0.000156999029337735
Rx227 x227 0 1
Fxc227_228 x227 0 Vx228 151.022608907286
Cx227 x227 xm227 1.0660761974355e-13
Vx227 xm227 0 0
Gx227_2 x227 0 u2 0 -7.37554054920054e-08
Rx228 x228 0 1
Fxc228_227 x228 0 Vx227 -411.070910718945
Cx228 x228 xm228 1.0660761974355e-13
Vx228 xm228 0 0
Gx228_2 x228 0 u2 0 3.03187017060438e-05
Rx229 x229 0 1
Fxc229_230 x229 0 Vx230 286.386072154125
Cx229 x229 xm229 6.29358278007233e-14
Vx229 xm229 0 0
Gx229_2 x229 0 u2 0 -1.52758721836916e-08
Rx230 x230 0 1
Fxc230_229 x230 0 Vx229 -652.184060451537
Cx230 x230 xm230 6.29358278007233e-14
Vx230 xm230 0 0
Gx230_2 x230 0 u2 0 9.96268034769865e-06
Rx231 x231 0 1
Fxc231_232 x231 0 Vx232 370.304622748678
Cx231 x231 xm231 6.18092938643569e-14
Vx231 xm231 0 0
Gx231_2 x231 0 u2 0 -1.80770398246959e-08
Rx232 x232 0 1
Fxc232_231 x232 0 Vx231 -546.029263057993
Cx232 x232 xm232 6.18092938643569e-14
Vx232 xm232 0 0
Gx232_2 x232 0 u2 0 9.87059273374871e-06
Rx233 x233 0 1
Fxc233_234 x233 0 Vx234 491.538446760153
Cx233 x233 xm233 5.92714932806977e-14
Vx233 xm233 0 0
Gx233_2 x233 0 u2 0 -2.42821917817464e-08
Rx234 x234 0 1
Fxc234_233 x234 0 Vx233 -467.056439549113
Cx234 x234 xm234 5.92714932806977e-14
Vx234 xm234 0 0
Gx234_2 x234 0 u2 0 1.13411540380312e-05
Rx235 x235 0 1
Fxc235_236 x235 0 Vx236 39.5355392557215
Cx235 x235 xm235 4.85449289847599e-13
Vx235 xm235 0 0
Gx235_2 x235 0 u2 0 -2.78073024394091e-06
Rx236 x236 0 1
Fxc236_235 x236 0 Vx235 -88.8000915937169
Cx236 x236 xm236 4.85449289847599e-13
Vx236 xm236 0 0
Gx236_2 x236 0 u2 0 0.000246929100359372
Rx237 x237 0 1
Fxc237_238 x237 0 Vx238 261.421097054904
Cx237 x237 xm237 7.07373676456137e-14
Vx237 xm237 0 0
Gx237_2 x237 0 u2 0 -1.71176773075854e-08
Rx238 x238 0 1
Fxc238_237 x238 0 Vx237 -630.769647347427
Cx238 x238 xm238 7.07373676456137e-14
Vx238 xm238 0 0
Gx238_2 x238 0 u2 0 1.07973112787127e-05
Rx239 x239 0 1
Fxc239_240 x239 0 Vx240 888.780289183778
Cx239 x239 xm239 4.92699889036898e-14
Vx239 xm239 0 0
Gx239_2 x239 0 u2 0 -1.87086836462519e-08
Rx240 x240 0 1
Fxc240_239 x240 0 Vx239 -400.718113932689
Cx240 x240 xm240 4.92699889036898e-14
Vx240 xm240 0 0
Gx240_2 x240 0 u2 0 7.49690842488941e-06
Rx241 x241 0 1
Fxc241_242 x241 0 Vx242 284.738363436963
Cx241 x241 xm241 1.55367016383078e-13
Vx241 xm241 0 0
Gx241_2 x241 0 u2 0 -1.12379520331441e-07
Rx242 x242 0 1
Fxc242_241 x242 0 Vx241 -130.135547688063
Cx242 x242 xm242 1.55367016383078e-13
Vx242 xm242 0 0
Gx242_2 x242 0 u2 0 1.4624570427254e-05
Rx243 x243 0 1
Fxc243_244 x243 0 Vx244 337.175946186913
Cx243 x243 xm243 8.2745464547176e-14
Vx243 xm243 0 0
Gx243_2 x243 0 u2 0 -2.64839285748991e-08
Rx244 x244 0 1
Fxc244_243 x244 0 Vx243 -403.983719929936
Cx244 x244 xm244 8.2745464547176e-14
Vx244 xm244 0 0
Gx244_2 x244 0 u2 0 1.06990759840465e-05
Rx245 x245 0 1
Fxc245_246 x245 0 Vx246 196.571273453853
Cx245 x245 xm245 1.78520263333676e-13
Vx245 xm245 0 0
Gx245_2 x245 0 u2 0 -2.29476109555537e-07
Rx246 x246 0 1
Fxc246_245 x246 0 Vx245 -153.37285659584
Cx246 x246 xm246 1.78520263333676e-13
Vx246 xm246 0 0
Gx246_2 x246 0 u2 0 3.51954064430327e-05
Rx247 x247 0 1
Fxc247_248 x247 0 Vx248 486.636880108467
Cx247 x247 xm247 1.06144284233908e-13
Vx247 xm247 0 0
Gx247_2 x247 0 u2 0 -5.08987852161311e-08
Rx248 x248 0 1
Fxc248_247 x248 0 Vx247 -178.223731563797
Cx248 x248 xm248 1.06144284233908e-13
Vx248 xm248 0 0
Gx248_2 x248 0 u2 0 9.07137143328313e-06
Rx249 x249 0 1
Fxc249_250 x249 0 Vx250 0.312174380362878
Cx249 x249 xm249 4.03773986408564e-11
Vx249 xm249 0 0
Gx249_2 x249 0 u2 0 -3.69444464968164
Rx250 x250 0 1
Fxc250_249 x250 0 Vx249 -0.642931026012734
Cx250 x250 xm250 4.03773986408564e-11
Vx250 xm250 0 0
Gx250_2 x250 0 u2 0 2.37527308916707
Rx251 x251 0 1
Fxc251_252 x251 0 Vx252 327.512364416066
Cx251 x251 xm251 4.28734109622567e-14
Vx251 xm251 0 0
Gx251_2 x251 0 u2 0 -4.21003556402675e-09
Rx252 x252 0 1
Fxc252_251 x252 0 Vx251 -1682.1829070575
Cx252 x252 xm252 4.28734109622567e-14
Vx252 xm252 0 0
Gx252_2 x252 0 u2 0 7.08204986390997e-06
Rx253 x253 0 1
Fxc253_254 x253 0 Vx254 431.532640274304
Cx253 x253 xm253 3.84734228551788e-14
Vx253 xm253 0 0
Gx253_2 x253 0 u2 0 -2.32255546122113e-09
Rx254 x254 0 1
Fxc254_253 x254 0 Vx253 -1654.83331130004
Cx254 x254 xm254 3.84734228551787e-14
Vx254 xm254 0 0
Gx254_2 x254 0 u2 0 3.84344214457056e-06
Rx255 x255 0 1
Fxc255_256 x255 0 Vx256 9.05713932066163
Cx255 x255 xm255 2.41483364210631e-12
Vx255 xm255 0 0
Gx255_2 x255 0 u2 0 -0.000165212259151167
Rx256 x256 0 1
Fxc256_255 x256 0 Vx255 -21.2964680553188
Cx256 x256 xm256 2.41483364210631e-12
Vx256 xm256 0 0
Gx256_2 x256 0 u2 0 0.00351843759935987
Rx257 x257 0 1
Fxc257_258 x257 0 Vx258 76.695620411658
Cx257 x257 xm257 3.4976618046498e-13
Vx257 xm257 0 0
Gx257_2 x257 0 u2 0 -4.20966582057393e-07
Rx258 x258 0 1
Fxc258_257 x258 0 Vx257 -117.135667459045
Cx258 x258 xm258 3.4976618046498e-13
Vx258 xm258 0 0
Gx258_2 x258 0 u2 0 4.93102015672454e-05
Rx259 x259 0 1
Fxc259_260 x259 0 Vx260 775.857623730808
Cx259 x259 xm259 1.82634891235488e-14
Vx259 xm259 0 0
Gx259_2 x259 0 u2 0 -4.92365148151007e-10
Rx260 x260 0 1
Fxc260_259 x260 0 Vx259 -4349.64211090205
Cx260 x260 xm260 1.82634891235488e-14
Vx260 xm260 0 0
Gx260_2 x260 0 u2 0 2.14161218233815e-06
Rx261 x261 0 1
Fxc261_262 x261 0 Vx262 2525.93067065548
Cx261 x261 xm261 8.73129447755975e-14
Vx261 xm261 0 0
Gx261_2 x261 0 u2 0 -3.27437506280311e-08
Rx262 x262 0 1
Fxc262_261 x262 0 Vx261 -60.9726961850079
Cx262 x262 xm262 8.73129447755975e-14
Vx262 xm262 0 0
Gx262_2 x262 0 u2 0 1.9964747590006e-06
Rx263 x263 0 1
Fxc263_264 x263 0 Vx264 9.73300514757486
Cx263 x263 xm263 1.19432876562705e-11
Vx263 xm263 0 0
Gx263_2 x263 0 u2 0 -0.0702844413961561
Rx264 x264 0 1
Fxc264_263 x264 0 Vx263 -1.12210195431616
Cx264 x264 xm264 1.19432876562705e-11
Vx264 xm264 0 0
Gx264_2 x264 0 u2 0 0.0788663090486463
Rx265 x265 0 1
Fxc265_266 x265 0 Vx266 126.623385780357
Cx265 x265 xm265 2.49726015690021e-13
Vx265 xm265 0 0
Gx265_2 x265 0 u2 0 -3.04798131315897e-07
Rx266 x266 0 1
Fxc266_265 x266 0 Vx265 -155.211672463462
Cx266 x266 xm266 2.49726015690021e-13
Vx266 xm266 0 0
Gx266_2 x266 0 u2 0 4.73082277252784e-05
Rx267 x267 0 1
Fxc267_268 x267 0 Vx268 1726.09143040798
Cx267 x267 xm267 2.53897718170844e-14
Vx267 xm267 0 0
Gx267_2 x267 0 u2 0 -1.38283911286938e-09
Rx268 x268 0 1
Fxc268_267 x268 0 Vx267 -1124.9686971473
Cx268 x268 xm268 2.53897718170844e-14
Vx268 xm268 0 0
Gx268_2 x268 0 u2 0 1.55565071516899e-06
Rx269 x269 0 1
Fxc269_270 x269 0 Vx270 0.830678964802864
Cx269 x269 xm269 2.12240440031949e-11
Vx269 xm269 0 0
Gx269_2 x269 0 u2 0 -0.18400999788669
Rx270 x270 0 1
Fxc270_269 x270 0 Vx269 -4.30416145879425
Cx270 x270 xm270 2.12240440031949e-11
Vx270 xm270 0 0
Gx270_2 x270 0 u2 0 0.792008740936703
Rx271 x271 0 1
Fxc271_272 x271 0 Vx272 366.153861842453
Cx271 x271 xm271 1.58125194797678e-13
Vx271 xm271 0 0
Gx271_2 x271 0 u2 0 -1.00709701507812e-07
Rx272 x272 0 1
Fxc272_271 x272 0 Vx271 -142.455629598624
Cx272 x272 xm272 1.58125194797678e-13
Vx272 xm272 0 0
Gx272_2 x272 0 u2 0 1.43466639349849e-05
Rx273 x273 0 1
Fxc273_274 x273 0 Vx274 212.535835986321
Cx273 x273 xm273 2.51123986719261e-13
Vx273 xm273 0 0
Gx273_2 x273 0 u2 0 -2.71268702997101e-07
Rx274 x274 0 1
Fxc274_273 x274 0 Vx273 -101.709668752464
Cx274 x274 xm274 2.51123986719261e-13
Vx274 xm274 0 0
Gx274_2 x274 0 u2 0 2.75906499247456e-05
Rx275 x275 0 1
Fxc275_276 x275 0 Vx276 1514.9682594056
Cx275 x275 xm275 5.50290062427746e-14
Vx275 xm275 0 0
Gx275_2 x275 0 u2 0 -5.24111165164938e-09
Rx276 x276 0 1
Fxc276_275 x276 0 Vx275 -305.086944063805
Cx276 x276 xm276 5.50290062427746e-14
Vx276 xm276 0 0
Gx276_2 x276 0 u2 0 1.59899473729891e-06
Rx277 x277 0 1
Fxc277_278 x277 0 Vx278 130.540989317584
Cx277 x277 xm277 1.73036537262631e-13
Vx277 xm277 0 0
Gx277_2 x277 0 u2 0 -6.49867431095607e-08
Rx278 x278 0 1
Fxc278_277 x278 0 Vx277 -372.881443758699
Cx278 x278 xm278 1.73036537262631e-13
Vx278 xm278 0 0
Gx278_2 x278 0 u2 0 2.42323505958687e-05
Rx279 x279 0 1
Fxc279_280 x279 0 Vx280 155.583209065286
Cx279 x279 xm279 1.04005943428604e-12
Vx279 xm279 0 0
Gx279_2 x279 0 u2 0 -1.18530059860113e-05
Rx280 x280 0 1
Fxc280_279 x280 0 Vx279 -8.86703180124089
Cx280 x280 xm280 1.04005943428604e-12
Vx280 xm280 0 0
Gx280_2 x280 0 u2 0 0.000105100981018261
Rx281 x281 0 1
Fxc281_282 x281 0 Vx282 164.485245709916
Cx281 x281 xm281 1.69597975933451e-13
Vx281 xm281 0 0
Gx281_2 x281 0 u2 0 -6.96509324215613e-08
Rx282 x282 0 1
Fxc282_281 x282 0 Vx281 -322.397763709952
Cx282 x282 xm282 1.69597975933451e-13
Vx282 xm282 0 0
Gx282_2 x282 0 u2 0 2.24553048530243e-05
Rx283 x283 0 1
Fxc283_284 x283 0 Vx284 198.975906585284
Cx283 x283 xm283 1.6574520023931e-13
Vx283 xm283 0 0
Gx283_2 x283 0 u2 0 -5.72183979893912e-08
Rx284 x284 0 1
Fxc284_283 x284 0 Vx283 -291.340814173171
Cx284 x284 xm284 1.6574520023931e-13
Vx284 xm284 0 0
Gx284_2 x284 0 u2 0 1.66700546559137e-05
Rx285 x285 0 1
Fxc285_286 x285 0 Vx286 608.30842567059
Cx285 x285 xm285 4.17930149743441e-14
Vx285 xm285 0 0
Gx285_2 x285 0 u2 0 -2.19000538189868e-09
Rx286 x286 0 1
Fxc286_285 x286 0 Vx285 -1572.1641490067
Cx286 x286 xm286 4.17930149743441e-14
Vx286 xm286 0 0
Gx286_2 x286 0 u2 0 3.44304794755283e-06
Rx287 x287 0 1
Fxc287_288 x287 0 Vx288 455.896506615464
Cx287 x287 xm287 9.47540753730688e-14
Vx287 xm287 0 0
Gx287_2 x287 0 u2 0 -1.6440864981683e-08
Rx288 x288 0 1
Fxc288_287 x288 0 Vx287 -420.361574203469
Cx288 x288 xm288 9.47540753730688e-14
Vx288 xm288 0 0
Gx288_2 x288 0 u2 0 6.91110788496694e-06
Rx289 x289 0 1
Fxc289_290 x289 0 Vx290 62.188749482855
Cx289 x289 xm289 3.39327012867075e-13
Vx289 xm289 0 0
Gx289_2 x289 0 u2 0 -1.2898790409243e-07
Rx290 x290 0 1
Fxc290_289 x290 0 Vx289 -248.752165049731
Cx290 x290 xm290 3.39327012867075e-13
Vx290 xm290 0 0
Gx290_2 x290 0 u2 0 3.20860204082191e-05
Rx291 x291 0 1
Fxc291_292 x291 0 Vx292 1483.73931434654
Cx291 x291 xm291 2.21690564685036e-14
Vx291 xm291 0 0
Gx291_2 x291 0 u2 0 -2.12674104529195e-09
Rx292 x292 0 1
Fxc292_291 x292 0 Vx291 -2511.44342893749
Cx292 x292 xm292 2.21690564685036e-14
Vx292 xm292 0 0
Gx292_2 x292 0 u2 0 5.34118982325012e-06
Rx293 x293 0 1
Fxc293_294 x293 0 Vx294 301.860036929104
Cx293 x293 xm293 1.4311943973241e-13
Vx293 xm293 0 0
Gx293_2 x293 0 u2 0 -2.49345234552723e-08
Rx294 x294 0 1
Fxc294_293 x294 0 Vx293 -312.403154879864
Cx294 x294 xm294 1.4311943973241e-13
Vx294 xm294 0 0
Gx294_2 x294 0 u2 0 7.78962379285304e-06
Rx295 x295 0 1
Fxc295_296 x295 0 Vx296 517.12127884219
Cx295 x295 xm295 1.49527034425067e-14
Vx295 xm295 0 0
Gx295_2 x295 0 u2 0 -7.55830037472335e-10
Rx296 x296 0 1
Fxc296_295 x296 0 Vx295 -17416.7527408689
Cx296 x296 xm296 1.49527034425067e-14
Vx296 xm296 0 0
Gx296_2 x296 0 u2 0 1.31641048767774e-05
Rx297 x297 0 1
Fxc297_298 x297 0 Vx298 257.876917626468
Cx297 x297 xm297 1.29249231176747e-13
Vx297 xm297 0 0
Gx297_2 x297 0 u2 0 -1.89467370341867e-08
Rx298 x298 0 1
Fxc298_297 x298 0 Vx297 -485.254097869213
Cx298 x298 xm298 1.29249231176747e-13
Vx298 xm298 0 0
Gx298_2 x298 0 u2 0 9.19398178708946e-06
Rx299 x299 0 1
Fxc299_300 x299 0 Vx300 326.960855263058
Cx299 x299 xm299 2.97577142965506e-14
Vx299 xm299 0 0
Gx299_2 x299 0 u2 0 -1.02477206260601e-09
Rx300 x300 0 1
Fxc300_299 x300 0 Vx299 -7494.66462789677
Cx300 x300 xm300 2.97577142965506e-14
Vx300 xm300 0 0
Gx300_2 x300 0 u2 0 7.68032292927005e-06
Rx301 x301 0 1
Fxc301_302 x301 0 Vx302 277.922161908866
Cx301 x301 xm301 3.66480875628994e-13
Vx301 xm301 0 0
Gx301_2 x301 0 u2 0 -2.58733732741993e-07
Rx302 x302 0 1
Fxc302_301 x302 0 Vx301 -60.2545018482701
Cx302 x302 xm302 3.66480875628994e-13
Vx302 xm302 0 0
Gx302_2 x302 0 u2 0 1.55898721777123e-05
Rx303 x303 0 1
Fxc303_304 x303 0 Vx304 342.505849593461
Cx303 x303 xm303 1.55725403798337e-13
Vx303 xm303 0 0
Gx303_2 x303 0 u2 0 -3.78871016531309e-08
Rx304 x304 0 1
Fxc304_303 x304 0 Vx303 -282.211781610062
Cx304 x304 xm304 1.55725403798336e-13
Vx304 xm304 0 0
Gx304_2 x304 0 u2 0 1.06921864575716e-05
Rx305 x305 0 1
Fxc305_306 x305 0 Vx306 2693.96267389885
Cx305 x305 xm305 2.70690945024366e-14
Vx305 xm305 0 0
Gx305_2 x305 0 u2 0 -4.31048748723009e-09
Rx306 x306 0 1
Fxc306_305 x306 0 Vx305 -1302.9965321441
Cx306 x306 xm306 2.70690945024366e-14
Vx306 xm306 0 0
Gx306_2 x306 0 u2 0 5.61655024771133e-06
Rx307 x307 0 1
Fxc307_308 x307 0 Vx308 436.916845005531
Cx307 x307 xm307 1.05947857159888e-13
Vx307 xm307 0 0
Gx307_2 x307 0 u2 0 -1.16083449272805e-08
Rx308 x308 0 1
Fxc308_307 x308 0 Vx307 -503.25527716541
Cx308 x308 xm308 1.05947857159888e-13
Vx308 xm308 0 0
Gx308_2 x308 0 u2 0 5.84196084381024e-06
Rx309 x309 0 1
Fxc309_310 x309 0 Vx310 488.43030877387
Cx309 x309 xm309 8.05411899100067e-14
Vx309 xm309 0 0
Gx309_2 x309 0 u2 0 -5.06821476301497e-09
Rx310 x310 0 1
Fxc310_309 x310 0 Vx309 -868.274542170374
Cx310 x310 xm310 8.05411899100067e-14
Vx310 xm310 0 0
Gx310_2 x310 0 u2 0 4.40060185297795e-06
Rx311 x311 0 1
Fxc311_312 x311 0 Vx312 390.989647807331
Cx311 x311 xm311 2.77463484357731e-13
Vx311 xm311 0 0
Gx311_2 x311 0 u2 0 -1.23788289456569e-07
Rx312 x312 0 1
Fxc312_311 x312 0 Vx311 -94.6558922303475
Cx312 x312 xm312 2.77463484357731e-13
Vx312 xm312 0 0
Gx312_2 x312 0 u2 0 1.17172909861801e-05
Rx313 x313 0 1
Cx313 x313 0 1.26327330229509e-10
Gx313_2 x313 0 u2 0 -0.897951049739533
Rx314 x314 0 1
Fxc314_315 x314 0 Vx315 210.901279882153
Cx314 x314 xm314 1.99280702854811e-13
Vx314 xm314 0 0
Gx314_2 x314 0 u2 0 -3.63644689261627e-08
Rx315 x315 0 1
Fxc315_314 x315 0 Vx314 -356.108361883805
Cx315 x315 xm315 1.99280702854811e-13
Vx315 xm315 0 0
Gx315_2 x315 0 u2 0 1.29496914600703e-05
Rx316 x316 0 1
Fxc316_317 x316 0 Vx317 1409.32725263913
Cx316 x316 xm316 3.34725367390173e-14
Vx316 xm316 0 0
Gx316_2 x316 0 u2 0 -4.74327580008424e-09
Rx317 x317 0 1
Fxc317_316 x317 0 Vx316 -1993.88094552994
Cx317 x317 xm317 3.34725367390173e-14
Vx317 xm317 0 0
Gx317_2 x317 0 u2 0 9.45752723718123e-06
Rx318 x318 0 1
Fxc318_319 x318 0 Vx319 49.4897241135416
Cx318 x318 xm318 1.20981905835219e-12
Vx318 xm318 0 0
Gx318_2 x318 0 u2 0 -2.41501378831431e-06
Rx319 x319 0 1
Fxc319_318 x319 0 Vx318 -44.9127280459785
Cx319 x319 xm319 1.20981905835219e-12
Vx319 xm319 0 0
Gx319_2 x319 0 u2 0 0.000108464857501849
Rx320 x320 0 1
Fxc320_321 x320 0 Vx321 269.43162426058
Cx320 x320 xm320 2.41747187333388e-13
Vx320 xm320 0 0
Gx320_2 x320 0 u2 0 -4.4973451703016e-08
Rx321 x321 0 1
Fxc321_320 x321 0 Vx320 -223.370436799713
Cx321 x321 xm321 2.41747187333388e-13
Vx321 xm321 0 0
Gx321_2 x321 0 u2 0 1.00457395512935e-05
Rx322 x322 0 1
Fxc322_323 x322 0 Vx323 84.6749962408462
Cx322 x322 xm322 6.05595987313277e-13
Vx322 xm322 0 0
Gx322_2 x322 0 u2 0 -3.80956835421622e-07
Rx323 x323 0 1
Fxc323_322 x323 0 Vx322 -115.835982759894
Cx323 x323 xm323 6.05595987313277e-13
Vx323 xm323 0 0
Gx323_2 x323 0 u2 0 4.41285094201627e-05
Rx324 x324 0 1
Fxc324_325 x324 0 Vx325 10.2985665105747
Cx324 x324 xm324 4.27273098109608e-12
Vx324 xm324 0 0
Gx324_2 x324 0 u2 0 -6.67907787224067e-05
Rx325 x325 0 1
Fxc325_324 x325 0 Vx324 -22.3608649639
Cx325 x325 xm325 4.27273098109608e-12
Vx325 xm325 0 0
Gx325_2 x325 0 u2 0 0.00149349958384546
Rx326 x326 0 1
Fxc326_327 x326 0 Vx327 300.187541412766
Cx326 x326 xm326 2.2113064440014e-13
Vx326 xm326 0 0
Gx326_2 x326 0 u2 0 -1.85972749382598e-08
Rx327 x327 0 1
Fxc327_326 x327 0 Vx326 -266.169475136405
Cx327 x327 xm327 2.2113064440014e-13
Vx327 xm327 0 0
Gx327_2 x327 0 u2 0 4.95002690928405e-06
Rx328 x328 0 1
Fxc328_329 x328 0 Vx329 182.250067961427
Cx328 x328 xm328 3.84635353963742e-13
Vx328 xm328 0 0
Gx328_2 x328 0 u2 0 -1.04997391299436e-07
Rx329 x329 0 1
Fxc329_328 x329 0 Vx328 -152.224864183209
Cx329 x329 xm329 3.84635353963742e-13
Vx329 xm329 0 0
Gx329_2 x329 0 u2 0 1.59832136301479e-05
Rx330 x330 0 1
Fxc330_331 x330 0 Vx331 27.5863711311736
Cx330 x330 xm330 1.31174697600352e-12
Vx330 xm330 0 0
Gx330_2 x330 0 u2 0 -3.79888920425862e-06
Rx331 x331 0 1
Fxc331_330 x331 0 Vx330 -91.889884776176
Cx331 x331 xm331 1.31174697600352e-12
Vx331 xm331 0 0
Gx331_2 x331 0 u2 0 0.000349079491256783
Rx332 x332 0 1
Fxc332_333 x332 0 Vx333 139.206597722383
Cx332 x332 xm332 6.73245820833979e-13
Vx332 xm332 0 0
Gx332_2 x332 0 u2 0 -8.89805849488631e-07
Rx333 x333 0 1
Fxc333_332 x333 0 Vx332 -70.345328431322
Cx333 x333 xm333 6.73245820833979e-13
Vx333 xm333 0 0
Gx333_2 x333 0 u2 0 6.25936847223892e-05
Rx334 x334 0 1
Fxc334_335 x334 0 Vx335 416.30188641895
Cx334 x334 xm334 5.84808784752663e-13
Vx334 xm334 0 0
Gx334_2 x334 0 u2 0 -2.05200798447006e-07
Rx335 x335 0 1
Fxc335_334 x335 0 Vx334 -34.3643808465372
Cx335 x335 xm335 5.84808784752663e-13
Vx335 xm335 0 0
Gx335_2 x335 0 u2 0 7.05159838784644e-06
Rx336 x336 0 1
Fxc336_337 x336 0 Vx337 247.195134583799
Cx336 x336 xm336 1.79416446898388e-13
Vx336 xm336 0 0
Gx336_2 x336 0 u2 0 -1.34610327019602e-08
Rx337 x337 0 1
Fxc337_336 x337 0 Vx336 -671.577917544577
Cx337 x337 xm337 1.79416446898388e-13
Vx337 xm337 0 0
Gx337_2 x337 0 u2 0 9.04013230998192e-06
Rx338 x338 0 1
Fxc338_339 x338 0 Vx339 158.62242692603
Cx338 x338 xm338 9.55321996041439e-13
Vx338 xm338 0 0
Gx338_2 x338 0 u2 0 -6.4944982769255e-07
Rx339 x339 0 1
Fxc339_338 x339 0 Vx338 -40.3337594204834
Cx339 x339 xm339 9.55321996041439e-13
Vx339 xm339 0 0
Gx339_2 x339 0 u2 0 2.61947531058258e-05
Rx340 x340 0 1
Fxc340_341 x340 0 Vx341 95.7101534317422
Cx340 x340 xm340 4.22656817502044e-13
Vx340 xm340 0 0
Gx340_2 x340 0 u2 0 -6.2188553919407e-08
Rx341 x341 0 1
Fxc341_340 x341 0 Vx340 -353.718066150987
Cx341 x341 xm341 4.22656817502044e-13
Vx341 xm341 0 0
Gx341_2 x341 0 u2 0 2.1997215029099e-05
Rx342 x342 0 1
Fxc342_343 x342 0 Vx343 66.147544741668
Cx342 x342 xm342 2.32688864615857e-12
Vx342 xm342 0 0
Gx342_2 x342 0 u2 0 -4.78328518804739e-06
Rx343 x343 0 1
Fxc343_342 x343 0 Vx342 -18.5179155981617
Cx343 x343 xm343 2.32688864615857e-12
Vx343 xm343 0 0
Gx343_2 x343 0 u2 0 8.85764713941983e-05
Rx344 x344 0 1
Fxc344_345 x344 0 Vx345 1744.21789783878
Cx344 x344 xm344 2.24826805546157e-13
Vx344 xm344 0 0
Gx344_2 x344 0 u2 0 -2.15031547608821e-08
Rx345 x345 0 1
Fxc345_344 x345 0 Vx344 -75.5555524389227
Cx345 x345 xm345 2.24826805546157e-13
Vx345 xm345 0 0
Gx345_2 x345 0 u2 0 1.6246827371381e-06
Rx346 x346 0 1
Fxc346_347 x346 0 Vx347 135.804315286581
Cx346 x346 xm346 7.62490228495289e-13
Vx346 xm346 0 0
Gx346_2 x346 0 u2 0 -1.95678145291133e-07
Rx347 x347 0 1
Fxc347_346 x347 0 Vx346 -95.5071419423708
Cx347 x347 xm347 7.62490228495289e-13
Vx347 xm347 0 0
Gx347_2 x347 0 u2 0 1.86886603973401e-05
Rx348 x348 0 1
Fxc348_349 x348 0 Vx349 82.0064077344706
Cx348 x348 xm348 3.12815339647046e-13
Vx348 xm348 0 0
Gx348_2 x348 0 u2 0 -9.70340725688157e-09
Rx349 x349 0 1
Fxc349_348 x349 0 Vx348 -1022.86623563955
Cx349 x349 xm349 3.12815339647046e-13
Vx349 xm349 0 0
Gx349_2 x349 0 u2 0 9.92528765372398e-06
Rx350 x350 0 1
Fxc350_351 x350 0 Vx351 34.7581074079482
Cx350 x350 xm350 1.21980473796757e-12
Vx350 xm350 0 0
Gx350_2 x350 0 u2 0 -1.98913065529147e-07
Rx351 x351 0 1
Fxc351_350 x351 0 Vx350 -166.649294041749
Cx351 x351 xm351 1.21980473796757e-12
Vx351 xm351 0 0
Gx351_2 x351 0 u2 0 3.31487219461125e-05
Rx352 x352 0 1
Fxc352_353 x352 0 Vx353 5.60226483340145
Cx352 x352 xm352 6.30927595670662e-12
Vx352 xm352 0 0
Gx352_2 x352 0 u2 0 -1.33654803744237e-05
Rx353 x353 0 1
Fxc353_352 x353 0 Vx352 -45.6884954688949
Cx353 x353 xm353 6.30927595670662e-12
Vx353 xm353 0 0
Gx353_2 x353 0 u2 0 0.00061064868952646
Rx354 x354 0 1
Fxc354_355 x354 0 Vx355 7264.38816971335
Cx354 x354 xm354 5.94898906330198e-14
Vx354 xm354 0 0
Gx354_2 x354 0 u2 0 -1.60755461465736e-08
Rx355 x355 0 1
Fxc355_354 x355 0 Vx354 -388.010874944369
Cx355 x355 xm355 5.94898906330198e-14
Vx355 xm355 0 0
Gx355_2 x355 0 u2 0 6.23748672554061e-06
Rx356 x356 0 1
Fxc356_357 x356 0 Vx357 83.8984878757303
Cx356 x356 xm356 1.88629779420802e-12
Vx356 xm356 0 0
Gx356_2 x356 0 u2 0 -1.11578257187626e-06
Rx357 x357 0 1
Fxc357_356 x357 0 Vx356 -36.5676864050964
Cx357 x357 xm357 1.88629779420802e-12
Vx357 xm357 0 0
Gx357_2 x357 0 u2 0 4.08015871846432e-05
Rx358 x358 0 1
Fxc358_359 x358 0 Vx359 32.4479134913414
Cx358 x358 xm358 2.53255697284169e-12
Vx358 xm358 0 0
Gx358_2 x358 0 u2 0 -1.67667897860464e-06
Rx359 x359 0 1
Fxc359_358 x359 0 Vx358 -61.7016805571644
Cx359 x359 xm359 2.53255697284169e-12
Vx359 xm359 0 0
Gx359_2 x359 0 u2 0 0.000103453910734776
Rx360 x360 0 1
Fxc360_361 x360 0 Vx361 39.6682507542863
Cx360 x360 xm360 1.07068178225324e-12
Vx360 xm360 0 0
Gx360_2 x360 0 u2 0 -1.18885103541375e-07
Rx361 x361 0 1
Fxc361_360 x361 0 Vx360 -301.88315627795
Cx361 x361 xm361 1.07068178225324e-12
Vx361 xm361 0 0
Gx361_2 x361 0 u2 0 3.58894102915012e-05
Rx362 x362 0 1
Cx362 x362 0 5.22190407222509e-10
Gx362_2 x362 0 u2 0 -0.216757193055407
Rx363 x363 0 1
Fxc363_364 x363 0 Vx364 125.109435709331
Cx363 x363 xm363 1.10121754249303e-12
Vx363 xm363 0 0
Gx363_2 x363 0 u2 0 -1.33668775638944e-07
Rx364 x364 0 1
Fxc364_363 x364 0 Vx363 -110.206121172888
Cx364 x364 xm364 1.10121754249303e-12
Vx364 xm364 0 0
Gx364_2 x364 0 u2 0 1.4731117285097e-05
Rx365 x365 0 1
Fxc365_366 x365 0 Vx366 77.3626208525846
Cx365 x365 xm365 1.3584005978461e-12
Vx365 xm365 0 0
Gx365_2 x365 0 u2 0 -1.92398556318053e-07
Rx366 x366 0 1
Fxc366_365 x366 0 Vx365 -133.840772225952
Cx366 x366 xm366 1.35840059784609e-12
Vx366 xm366 0 0
Gx366_2 x366 0 u2 0 2.57507713527666e-05
Rx367 x367 0 1
Fxc367_368 x367 0 Vx368 2.7030076796841
Cx367 x367 xm367 1.37582820475616e-11
Vx367 xm367 0 0
Gx367_2 x367 0 u2 0 -1.66220494157343e-05
Rx368 x368 0 1
Fxc368_367 x368 0 Vx367 -51.593569674104
Cx368 x368 xm368 1.37582820475616e-11
Vx368 xm368 0 0
Gx368_2 x368 0 u2 0 0.000857590864657089
Rx369 x369 0 1
Fxc369_370 x369 0 Vx370 11.5244685328862
Cx369 x369 xm369 2.55525080407755e-12
Vx369 xm369 0 0
Gx369_2 x369 0 u2 0 -6.17296672275501e-07
Rx370 x370 0 1
Fxc370_369 x370 0 Vx369 -193.652910821066
Cx370 x370 xm370 2.55525080407755e-12
Vx370 xm370 0 0
Gx370_2 x370 0 u2 0 0.000119541297426308
Rx371 x371 0 1
Fxc371_372 x371 0 Vx372 12.2954608891883
Cx371 x371 xm371 3.52048110577458e-12
Vx371 xm371 0 0
Gx371_2 x371 0 u2 0 -6.2690537300025e-07
Rx372 x372 0 1
Fxc372_371 x372 0 Vx371 -143.576692089056
Cx372 x372 xm372 3.52048110577458e-12
Vx372 xm372 0 0
Gx372_2 x372 0 u2 0 9.0008999708232e-05
Rx373 x373 0 1
Fxc373_374 x373 0 Vx374 3.98146511744896
Cx373 x373 xm373 8.01925764208566e-11
Vx373 xm373 0 0
Gx373_2 x373 0 u2 0 -0.00544582178681248
Rx374 x374 0 1
Fxc374_373 x374 0 Vx373 -1.96187055913106
Cx374 x374 xm374 8.01925764208566e-11
Vx374 xm374 0 0
Gx374_2 x374 0 u2 0 0.0106839974338219
Rx375 x375 0 1
Fxc375_376 x375 0 Vx376 45.963668867458
Cx375 x375 xm375 1.34818539204243e-12
Vx375 xm375 0 0
Gx375_2 x375 0 u2 0 -7.01685755437572e-08
Rx376 x376 0 1
Fxc376_375 x376 0 Vx375 -328.343561993825
Cx376 x376 xm376 1.34818539204243e-12
Vx376 xm376 0 0
Gx376_2 x376 0 u2 0 2.30394000340701e-05
Rx377 x377 0 1
Fxc377_378 x377 0 Vx378 0.739478880582497
Cx377 x377 xm377 2.60286578934868e-10
Vx377 xm377 0 0
Gx377_2 x377 0 u2 0 -0.00870069344906375
Rx378 x378 0 1
Fxc378_377 x378 0 Vx377 -3.98060212059004
Cx378 x378 xm378 2.60286578934868e-10
Vx378 xm378 0 0
Gx378_2 x378 0 u2 0 0.034633998793947
Rx379 x379 0 1
Fxc379_380 x379 0 Vx380 20.7303613861312
Cx379 x379 xm379 1.94992797826926e-12
Vx379 xm379 0 0
Gx379_2 x379 0 u2 0 -5.76472289232728e-08
Rx380 x380 0 1
Fxc380_379 x380 0 Vx379 -434.355408225064
Cx380 x380 xm380 1.94992797826926e-12
Vx380 xm380 0 0
Gx380_2 x380 0 u2 0 2.50393856520119e-05
Rx381 x381 0 1
Fxc381_382 x381 0 Vx382 58.7969588177801
Cx381 x381 xm381 2.33413529363335e-12
Vx381 xm381 0 0
Gx381_2 x381 0 u2 0 -5.93056415754385e-08
Rx382 x382 0 1
Fxc382_381 x382 0 Vx381 -277.66831672903
Cx382 x382 xm382 2.33413529363335e-12
Vx382 xm382 0 0
Gx382_2 x382 0 u2 0 1.64672976687872e-05
Rx383 x383 0 1
Fxc383_384 x383 0 Vx384 23.6780769523624
Cx383 x383 xm383 1.72271737747677e-11
Vx383 xm383 0 0
Gx383_2 x383 0 u2 0 -2.92443525860546e-05
Rx384 x384 0 1
Fxc384_383 x384 0 Vx383 -8.79997892359445
Cx384 x384 xm384 1.72271737747677e-11
Vx384 xm384 0 0
Gx384_2 x384 0 u2 0 0.000257349686391445
Rx385 x385 0 1
Fxc385_386 x385 0 Vx386 106.947850719343
Cx385 x385 xm385 3.38373728470339e-12
Vx385 xm385 0 0
Gx385_2 x385 0 u2 0 -7.19649993515706e-07
Rx386 x386 0 1
Fxc386_385 x386 0 Vx385 -34.8068561117889
Cx386 x386 xm386 3.38373728470339e-12
Vx386 xm386 0 0
Gx386_2 x386 0 u2 0 2.5048753775151e-05
Rx387 x387 0 1
Fxc387_388 x387 0 Vx388 21.5465242525573
Cx387 x387 xm387 5.83456226648167e-12
Vx387 xm387 0 0
Gx387_2 x387 0 u2 0 -1.83145373986134e-07
Rx388 x388 0 1
Fxc388_387 x388 0 Vx387 -198.159389307524
Cx388 x388 xm388 5.83456226648167e-12
Vx388 xm388 0 0
Gx388_2 x388 0 u2 0 3.62919754635905e-05
Rx389 x389 0 1
Fxc389_390 x389 0 Vx390 57.300533413887
Cx389 x389 xm389 3.71913677806581e-11
Vx389 xm389 0 0
Gx389_2 x389 0 u2 0 -0.000535390646430594
Rx390 x390 0 1
Fxc390_389 x390 0 Vx389 -3.30357297896837
Cx390 x390 xm390 3.71913677806581e-11
Vx390 xm390 0 0
Gx390_2 x390 0 u2 0 0.00176870207274052
Rx391 x391 0 1
Fxc391_392 x391 0 Vx392 63.1913626294967
Cx391 x391 xm391 3.43647746350443e-11
Vx391 xm391 0 0
Gx391_2 x391 0 u2 0 -0.000428169899686359
Rx392 x392 0 1
Fxc392_391 x392 0 Vx391 -3.49133447050937
Cx392 x392 xm392 3.43647746350443e-11
Vx392 xm392 0 0
Gx392_2 x392 0 u2 0 0.00149488433000953
Rx393 x393 0 1
Fxc393_394 x393 0 Vx394 0.503713378327978
Cx393 x393 xm393 1.92407202503742e-10
Vx393 xm393 0 0
Gx393_2 x393 0 u2 0 -3.14308373836539e-05
Rx394 x394 0 1
Fxc394_393 x394 0 Vx393 -48.6717930694524
Cx394 x394 xm394 1.92407202503742e-10
Vx394 xm394 0 0
Gx394_2 x394 0 u2 0 0.00152979521313681
Rx395 x395 0 1
Fxc395_396 x395 0 Vx396 784.684854400283
Cx395 x395 xm395 8.89563374249556e-13
Vx395 xm395 0 0
Gx395_2 x395 0 u2 0 -7.72444643005713e-08
Rx396 x396 0 1
Fxc396_395 x396 0 Vx395 -95.0115478991752
Cx396 x396 xm396 8.89563374249556e-13
Vx396 xm396 0 0
Gx396_2 x396 0 u2 0 7.33911611983986e-06
Rx397 x397 0 1
Fxc397_398 x397 0 Vx398 3.66502476950047
Cx397 x397 xm397 1.38719414317867e-09
Vx397 xm397 0 0
Gx397_2 x397 0 u2 0 -0.030642919065343
Rx398 x398 0 1
Fxc398_397 x398 0 Vx397 -0.158940480356061
Cx398 x398 xm398 1.38719414317867e-09
Vx398 xm398 0 0
Gx398_2 x398 0 u2 0 0.00487040027575752
Rx399 x399 0 1
Cx399 x399 0 4.58826427740312e-07
Gx399_2 x399 0 u2 0 -0.642318793742956
Rx400 x400 0 1
Cx400 x400 0 7.53723517430562e-08
Gx400_2 x400 0 u2 0 -0.272469801350741
Rx401 x401 0 1
Fxc401_402 x401 0 Vx402 1.53532509240335
Cx401 x401 xm401 4.30686999129145e-12
Vx401 xm401 0 0
Gx401_3 x401 0 u3 0 -0.326670507913715
Rx402 x402 0 1
Fxc402_401 x402 0 Vx401 -10.9580431829534
Cx402 x402 xm402 4.30686999129145e-12
Vx402 xm402 0 0
Gx402_3 x402 0 u3 0 3.57966953231582
Rx403 x403 0 1
Fxc403_404 x403 0 Vx404 1.05716032943846
Cx403 x403 xm403 8.05342537957096e-12
Vx403 xm403 0 0
Gx403_3 x403 0 u3 0 -0.468039169088175
Rx404 x404 0 1
Fxc404_403 x404 0 Vx403 -8.13697776579889
Cx404 x404 xm404 8.05342537957096e-12
Vx404 xm404 0 0
Gx404_3 x404 0 u3 0 3.80842431239346
Rx405 x405 0 1
Fxc405_406 x405 0 Vx406 934.212247445619
Cx405 x405 xm405 2.88356300968449e-14
Vx405 xm405 0 0
Gx405_3 x405 0 u3 0 -6.35307971841051e-08
Rx406 x406 0 1
Fxc406_405 x406 0 Vx405 -685.161248282117
Cx406 x406 xm406 2.88356300968449e-14
Vx406 xm406 0 0
Gx406_3 x406 0 u3 0 4.35288403030195e-05
Rx407 x407 0 1
Fxc407_408 x407 0 Vx408 1110.88474194833
Cx407 x407 xm407 3.27807622205493e-15
Vx407 xm407 0 0
Gx407_3 x407 0 u3 0 -2.09338974781689e-10
Rx408 x408 0 1
Fxc408_407 x408 0 Vx407 -46263.6792398485
Cx408 x408 xm408 3.27807622205493e-15
Vx408 xm408 0 0
Gx408_3 x408 0 u3 0 9.68479118169879e-06
Rx409 x409 0 1
Fxc409_410 x409 0 Vx410 1114.69197141555
Cx409 x409 xm409 8.61037113698984e-14
Vx409 xm409 0 0
Gx409_3 x409 0 u3 0 -5.5027395054669e-07
Rx410 x410 0 1
Fxc410_409 x410 0 Vx409 -68.321211127136
Cx410 x410 xm410 8.61037113698984e-14
Vx410 xm410 0 0
Gx410_3 x410 0 u3 0 3.75953827530636e-05
Rx411 x411 0 1
Fxc411_412 x411 0 Vx412 250.300015292538
Cx411 x411 xm411 7.36385701297364e-14
Vx411 xm411 0 0
Gx411_3 x411 0 u3 0 -2.3201810588944e-07
Rx412 x412 0 1
Fxc412_411 x412 0 Vx411 -423.032736012222
Cx412 x412 xm412 7.36385701297364e-14
Vx412 xm412 0 0
Gx412_3 x412 0 u3 0 9.81512541387831e-05
Rx413 x413 0 1
Fxc413_414 x413 0 Vx414 2952.78723245788
Cx413 x413 xm413 2.83512527353486e-14
Vx413 xm413 0 0
Gx413_3 x413 0 u3 0 -3.65013119643172e-08
Rx414 x414 0 1
Fxc414_413 x414 0 Vx413 -250.543340093902
Cx414 x414 xm414 2.83512527353486e-14
Vx414 xm414 0 0
Gx414_3 x414 0 u3 0 9.14516061734952e-06
Rx415 x415 0 1
Fxc415_416 x415 0 Vx416 7.49287809924968
Cx415 x415 xm415 2.47015112633796e-12
Vx415 xm415 0 0
Gx415_3 x415 0 u3 0 -0.00655357447820783
Rx416 x416 0 1
Fxc416_415 x416 0 Vx415 -15.038874252522
Cx416 x416 xm416 2.47015112633796e-12
Vx416 xm416 0 0
Gx416_3 x416 0 u3 0 0.0985583824823048
Rx417 x417 0 1
Fxc417_418 x417 0 Vx418 55.664243432534
Cx417 x417 xm417 6.21082676967847e-14
Vx417 xm417 0 0
Gx417_3 x417 0 u3 0 -2.40968149627136e-08
Rx418 x418 0 1
Fxc418_417 x418 0 Vx417 -2873.67941692104
Cx418 x418 xm418 6.21082676967847e-14
Vx418 xm418 0 0
Gx418_3 x418 0 u3 0 6.92465211717052e-05
Rx419 x419 0 1
Fxc419_420 x419 0 Vx420 494.786304494797
Cx419 x419 xm419 6.88618151548846e-14
Vx419 xm419 0 0
Gx419_3 x419 0 u3 0 -1.53670961578925e-07
Rx420 x420 0 1
Fxc420_419 x420 0 Vx419 -273.06588650051
Cx420 x420 xm420 6.88618151548846e-14
Vx420 xm420 0 0
Gx420_3 x420 0 u3 0 4.19622973529348e-05
Rx421 x421 0 1
Fxc421_422 x421 0 Vx422 18130.1682584514
Cx421 x421 xm421 5.46774161318971e-15
Vx421 xm421 0 0
Gx421_3 x421 0 u3 0 -1.51457107660153e-09
Rx422 x422 0 1
Fxc422_421 x422 0 Vx421 -1207.15215381898
Cx422 x422 xm422 5.46774161318971e-15
Vx422 xm422 0 0
Gx422_3 x422 0 u3 0 1.82831773723146e-06
Rx423 x423 0 1
Fxc423_424 x423 0 Vx424 158.767974475016
Cx423 x423 xm423 1.19014549350492e-13
Vx423 xm423 0 0
Gx423_3 x423 0 u3 0 -3.83814742610781e-07
Rx424 x424 0 1
Fxc424_423 x424 0 Vx423 -298.343857718692
Cx424 x424 xm424 1.19014549350492e-13
Vx424 xm424 0 0
Gx424_3 x424 0 u3 0 0.000114508770959807
Rx425 x425 0 1
Fxc425_426 x425 0 Vx426 60.6802830560271
Cx425 x425 xm425 3.39580797038266e-13
Vx425 xm425 0 0
Gx425_3 x425 0 u3 0 -7.70502383969245e-06
Rx426 x426 0 1
Fxc426_425 x426 0 Vx425 -99.6479914045633
Cx426 x426 xm426 3.39580797038266e-13
Vx426 xm426 0 0
Gx426_3 x426 0 u3 0 0.000767790149349628
Rx427 x427 0 1
Fxc427_428 x427 0 Vx428 101.247445630551
Cx427 x427 xm427 1.0660761974355e-13
Vx427 xm427 0 0
Gx427_3 x427 0 u3 0 -1.92109188154514e-07
Rx428 x428 0 1
Fxc428_427 x428 0 Vx427 -613.161161706743
Cx428 x428 xm428 1.0660761974355e-13
Vx428 xm428 0 0
Gx428_3 x428 0 u3 0 0.000117793892983361
Rx429 x429 0 1
Fxc429_430 x429 0 Vx430 90.7410767688417
Cx429 x429 xm429 6.29358278007233e-14
Vx429 xm429 0 0
Gx429_3 x429 0 u3 0 -1.83321054744926e-08
Rx430 x430 0 1
Fxc430_429 x430 0 Vx429 -2058.34488684819
Cx430 x430 xm430 6.29358278007233e-14
Vx430 xm430 0 0
Gx430_3 x430 0 u3 0 3.77337955685835e-05
Rx431 x431 0 1
Fxc431_432 x431 0 Vx432 947.894629534713
Cx431 x431 xm431 6.18092938643569e-14
Vx431 xm431 0 0
Gx431_3 x431 0 u3 0 -8.15271189362913e-08
Rx432 x432 0 1
Fxc432_431 x432 0 Vx431 -213.311853413158
Cx432 x432 xm432 6.18092938643569e-14
Vx432 xm432 0 0
Gx432_3 x432 0 u3 0 1.73907008437353e-05
Rx433 x433 0 1
Fxc433_434 x433 0 Vx434 643.981280080351
Cx433 x433 xm433 5.92714932806977e-14
Vx433 xm433 0 0
Gx433_3 x433 0 u3 0 -6.83411286917917e-08
Rx434 x434 0 1
Fxc434_433 x434 0 Vx433 -356.495140381493
Cx434 x434 xm434 5.92714932806977e-14
Vx434 xm434 0 0
Gx434_3 x434 0 u3 0 2.43632802668099e-05
Rx435 x435 0 1
Fxc435_436 x435 0 Vx436 27.4044468403675
Cx435 x435 xm435 4.85449289847599e-13
Vx435 xm435 0 0
Gx435_3 x435 0 u3 0 -7.37384861903198e-06
Rx436 x436 0 1
Fxc436_435 x436 0 Vx435 -128.109117748861
Cx436 x436 xm436 4.85449289847599e-13
Vx436 xm436 0 0
Gx436_3 x436 0 u3 0 0.000944657240997847
Rx437 x437 0 1
Fxc437_438 x437 0 Vx438 452.01376463838
Cx437 x437 xm437 7.07373676456137e-14
Vx437 xm437 0 0
Gx437_3 x437 0 u3 0 -8.90928717265891e-08
Rx438 x438 0 1
Fxc438_437 x438 0 Vx437 -364.804141153577
Cx438 x438 xm438 7.07373676456137e-14
Vx438 xm438 0 0
Gx438_3 x438 0 u3 0 3.25014485531241e-05
Rx439 x439 0 1
Fxc439_440 x439 0 Vx440 368.358116085704
Cx439 x439 xm439 4.92699889036898e-14
Vx439 xm439 0 0
Gx439_3 x439 0 u3 0 -2.58284180283086e-08
Rx440 x440 0 1
Fxc440_439 x440 0 Vx439 -966.859003859737
Cx440 x440 xm440 4.92699889036898e-14
Vx440 xm440 0 0
Gx440_3 x440 0 u3 0 2.49724385261233e-05
Rx441 x441 0 1
Fxc441_442 x441 0 Vx442 79.2527210607939
Cx441 x441 xm441 1.55367016383078e-13
Vx441 xm441 0 0
Gx441_3 x441 0 u3 0 -1.86561779383387e-07
Rx442 x442 0 1
Fxc442_441 x442 0 Vx441 -467.549661105615
Cx442 x442 xm442 1.55367016383078e-13
Vx442 xm442 0 0
Gx442_3 x442 0 u3 0 8.72268967259633e-05
Rx443 x443 0 1
Fxc443_444 x443 0 Vx444 893.933559364587
Cx443 x443 xm443 8.2745464547176e-14
Vx443 xm443 0 0
Gx443_3 x443 0 u3 0 -8.46327778142531e-08
Rx444 x444 0 1
Fxc444_443 x444 0 Vx443 -152.375522302023
Cx444 x444 xm444 8.2745464547176e-14
Vx444 xm444 0 0
Gx444_3 x444 0 u3 0 1.28959637233178e-05
Rx445 x445 0 1
Fxc445_446 x445 0 Vx446 226.896253049889
Cx445 x445 xm445 1.78520263333676e-13
Vx445 xm445 0 0
Gx445_3 x445 0 u3 0 -7.0609451794601e-07
Rx446 x446 0 1
Fxc446_445 x446 0 Vx445 -132.874374649415
Cx446 x446 xm446 1.78520263333676e-13
Vx446 xm446 0 0
Gx446_3 x446 0 u3 0 9.38218675154562e-05
Rx447 x447 0 1
Fxc447_448 x447 0 Vx448 598.806642937229
Cx447 x447 xm447 1.06144284233908e-13
Vx447 xm447 0 0
Gx447_3 x447 0 u3 0 -1.89336553970807e-07
Rx448 x448 0 1
Fxc448_447 x448 0 Vx447 -144.838474510021
Cx448 x448 xm448 1.06144284233908e-13
Vx448 xm448 0 0
Gx448_3 x448 0 u3 0 2.7423217646116e-05
Rx449 x449 0 1
Fxc449_450 x449 0 Vx450 0.498814700465461
Cx449 x449 xm449 4.03773986408564e-11
Vx449 xm449 0 0
Gx449_3 x449 0 u3 0 -21.8117329577295
Rx450 x450 0 1
Fxc450_449 x450 0 Vx449 -0.402367040254244
Cx450 x450 xm450 4.03773986408564e-11
Vx450 xm450 0 0
Gx450_3 x450 0 u3 0 8.77632243301758
Rx451 x451 0 1
Fxc451_452 x451 0 Vx452 120.182547219409
Cx451 x451 xm451 4.28734109622567e-14
Vx451 xm451 0 0
Gx451_3 x451 0 u3 0 -3.59732647400105e-09
Rx452 x452 0 1
Fxc452_451 x452 0 Vx451 -4584.15730085073
Cx452 x452 xm452 4.28734109622567e-14
Vx452 xm452 0 0
Gx452_3 x452 0 u3 0 1.64907104193355e-05
Rx453 x453 0 1
Fxc453_454 x453 0 Vx454 5280.69672382562
Cx453 x453 xm453 3.84734228551787e-14
Vx453 xm453 0 0
Gx453_3 x453 0 u3 0 -1.9031999894623e-08
Rx454 x454 0 1
Fxc454_453 x454 0 Vx453 -135.231130547076
Cx454 x454 xm454 3.84734228551787e-14
Vx454 xm454 0 0
Gx454_3 x454 0 u3 0 2.57371886232169e-06
Rx455 x455 0 1
Fxc455_456 x455 0 Vx456 2.26638095346044
Cx455 x455 xm455 2.41483364210631e-12
Vx455 xm455 0 0
Gx455_3 x455 0 u3 0 -0.000159538119688587
Rx456 x456 0 1
Fxc456_455 x456 0 Vx455 -85.107085779438
Cx456 x456 xm456 2.41483364210631e-12
Vx456 xm456 0 0
Gx456_3 x456 0 u3 0 0.0135778244374268
Rx457 x457 0 1
Fxc457_458 x457 0 Vx458 191.164621091096
Cx457 x457 xm457 3.4976618046498e-13
Vx457 xm457 0 0
Gx457_3 x457 0 u3 0 -2.17597449097653e-06
Rx458 x458 0 1
Fxc458_457 x458 0 Vx457 -46.9950592156067
Cx458 x458 xm458 3.4976618046498e-13
Vx458 xm458 0 0
Gx458_3 x458 0 u3 0 0.000102260050055091
Rx459 x459 0 1
Fxc459_460 x459 0 Vx460 2130.28092822623
Cx459 x459 xm459 1.82634891235488e-14
Vx459 xm459 0 0
Gx459_3 x459 0 u3 0 -8.86240703700182e-10
Rx460 x460 0 1
Fxc460_459 x460 0 Vx459 -1584.15866542722
Cx460 x460 xm460 1.82634891235488e-14
Vx460 xm460 0 0
Gx460_3 x460 0 u3 0 1.40394589042096e-06
Rx461 x461 0 1
Fxc461_462 x461 0 Vx462 275.470502128894
Cx461 x461 xm461 8.73129447755975e-14
Vx461 xm461 0 0
Gx461_3 x461 0 u3 0 -4.02216054917178e-08
Rx462 x462 0 1
Fxc462_461 x462 0 Vx461 -559.090001201676
Cx462 x462 xm462 8.73129447755975e-14
Vx462 xm462 0 0
Gx462_3 x462 0 u3 0 2.24874974626978e-05
Rx463 x463 0 1
Fxc463_464 x463 0 Vx464 38.7245027337495
Cx463 x463 xm463 1.19432876562705e-11
Vx463 xm463 0 0
Gx463_3 x463 0 u3 0 -0.25766773489269
Rx464 x464 0 1
Fxc464_463 x464 0 Vx463 -0.282028775748349
Cx464 x464 xm464 1.19432876562705e-11
Vx464 xm464 0 0
Gx464_3 x464 0 u3 0 0.0726697158216356
Rx465 x465 0 1
Fxc465_466 x465 0 Vx466 309.026510273391
Cx465 x465 xm465 2.49726015690021e-13
Vx465 xm465 0 0
Gx465_3 x465 0 u3 0 -6.13037104674916e-07
Rx466 x466 0 1
Fxc466_465 x466 0 Vx465 -63.597868877231
Cx466 x466 xm466 2.49726015690021e-13
Vx466 xm466 0 0
Gx466_3 x466 0 u3 0 3.89878533999926e-05
Rx467 x467 0 1
Fxc467_468 x467 0 Vx468 3953.66081663791
Cx467 x467 xm467 2.53897718170844e-14
Vx467 xm467 0 0
Gx467_3 x467 0 u3 0 -7.3978984320771e-09
Rx468 x468 0 1
Fxc468_467 x468 0 Vx467 -491.139457247228
Cx468 x468 xm468 2.53897718170844e-14
Vx468 xm468 0 0
Gx468_3 x468 0 u3 0 3.63339982070047e-06
Rx469 x469 0 1
Fxc469_470 x469 0 Vx470 0.300227401536388
Cx469 x469 xm469 2.12240440031949e-11
Vx469 xm469 0 0
Gx469_3 x469 0 u3 0 -0.332531287180552
Rx470 x470 0 1
Fxc470_469 x470 0 Vx469 -11.9088942802653
Cx470 x470 xm470 2.12240440031949e-11
Vx470 xm470 0 0
Gx470_3 x470 0 u3 0 3.96007994391372
Rx471 x471 0 1
Fxc471_472 x471 0 Vx472 178.892004802741
Cx471 x471 xm471 1.58125194797678e-13
Vx471 xm471 0 0
Gx471_3 x471 0 u3 0 -1.21300255400084e-07
Rx472 x472 0 1
Fxc472_471 x472 0 Vx471 -291.576356228164
Cx472 x472 xm472 1.58125194797678e-13
Vx472 xm472 0 0
Gx472_3 x472 0 u3 0 3.53682864791021e-05
Rx473 x473 0 1
Fxc473_474 x473 0 Vx474 1243.24202384221
Cx473 x473 xm473 2.51123986719261e-13
Vx473 xm473 0 0
Gx473_3 x473 0 u3 0 -6.45631750040072e-07
Rx474 x474 0 1
Fxc474_473 x474 0 Vx473 -17.387563371925
Cx474 x474 xm474 2.51123986719261e-13
Vx474 xm474 0 0
Gx474_3 x474 0 u3 0 1.12259629687486e-05
Rx475 x475 0 1
Fxc475_476 x475 0 Vx476 2661.2965852714
Cx475 x475 xm475 5.50290062427746e-14
Vx475 xm475 0 0
Gx475_3 x475 0 u3 0 -2.03618679366496e-08
Rx476 x476 0 1
Fxc476_475 x476 0 Vx475 -173.673629302982
Cx476 x476 xm476 5.50290062427746e-14
Vx476 xm476 0 0
Gx476_3 x476 0 u3 0 3.53631950394596e-06
Rx477 x477 0 1
Fxc477_478 x477 0 Vx478 162.837431846778
Cx477 x477 xm477 1.73036537262631e-13
Vx477 xm477 0 0
Gx477_3 x477 0 u3 0 -1.61605891476766e-07
Rx478 x478 0 1
Fxc478_477 x478 0 Vx477 -298.925818310817
Cx478 x478 xm478 1.73036537262631e-13
Vx478 xm478 0 0
Gx478_3 x478 0 u3 0 4.83081733535414e-05
Rx479 x479 0 1
Fxc479_480 x479 0 Vx480 161.039460670871
Cx479 x479 xm479 1.04005943428604e-12
Vx479 xm479 0 0
Gx479_3 x479 0 u3 0 -3.3166672601175e-05
Rx480 x480 0 1
Fxc480_479 x480 0 Vx479 -8.56660384215098
Cx480 x480 xm480 1.04005943428604e-12
Vx480 xm480 0 0
Gx480_3 x480 0 u3 0 0.00028412574493659
Rx481 x481 0 1
Fxc481_482 x481 0 Vx482 198.080229568018
Cx481 x481 xm481 1.69597975933452e-13
Vx481 xm481 0 0
Gx481_3 x481 0 u3 0 -1.52973576094286e-07
Rx482 x482 0 1
Fxc482_481 x482 0 Vx481 -267.718163977335
Cx482 x482 xm482 1.69597975933452e-13
Vx482 xm482 0 0
Gx482_3 x482 0 u3 0 4.09538049290093e-05
Rx483 x483 0 1
Fxc483_484 x483 0 Vx484 502.972779870991
Cx483 x483 xm483 1.6574520023931e-13
Vx483 xm483 0 0
Gx483_3 x483 0 u3 0 -1.16541594774536e-07
Rx484 x484 0 1
Fxc484_483 x484 0 Vx483 -115.254353605915
Cx484 x484 xm484 1.6574520023931e-13
Vx484 xm484 0 0
Gx484_3 x484 0 u3 0 1.34319261739417e-05
Rx485 x485 0 1
Fxc485_486 x485 0 Vx486 473.120171873981
Cx485 x485 xm485 4.17930149743441e-14
Vx485 xm485 0 0
Gx485_3 x485 0 u3 0 -4.3103968772076e-09
Rx486 x486 0 1
Fxc486_485 x486 0 Vx485 -2021.39066400395
Cx486 x486 xm486 4.17930149743441e-14
Vx486 xm486 0 0
Gx486_3 x486 0 u3 0 8.71299600573922e-06
Rx487 x487 0 1
Fxc487_488 x487 0 Vx488 342.431200394658
Cx487 x487 xm487 9.47540753730688e-14
Vx487 xm487 0 0
Gx487_3 x487 0 u3 0 -2.18097153969779e-08
Rx488 x488 0 1
Fxc488_487 x488 0 Vx487 -559.649275456993
Cx488 x488 xm488 9.47540753730688e-14
Vx488 xm488 0 0
Gx488_3 x488 0 u3 0 1.22057914198419e-05
Rx489 x489 0 1
Fxc489_490 x489 0 Vx490 55.4273555070049
Cx489 x489 xm489 3.39327012867075e-13
Vx489 xm489 0 0
Gx489_3 x489 0 u3 0 -2.79197744901999e-07
Rx490 x490 0 1
Fxc490_489 x490 0 Vx489 -279.096592902407
Cx490 x490 xm490 3.39327012867075e-13
Vx490 xm490 0 0
Gx490_3 x490 0 u3 0 7.79231393481833e-05
Rx491 x491 0 1
Fxc491_492 x491 0 Vx492 919.94133304292
Cx491 x491 xm491 2.21690564685036e-14
Vx491 xm491 0 0
Gx491_3 x491 0 u3 0 -2.83580418312048e-09
Rx492 x492 0 1
Fxc492_491 x492 0 Vx491 -4050.61411790918
Cx492 x492 xm492 2.21690564685036e-14
Vx492 xm492 0 0
Gx492_3 x492 0 u3 0 1.14867484597737e-05
Rx493 x493 0 1
Fxc493_494 x493 0 Vx494 675.394619132651
Cx493 x493 xm493 1.4311943973241e-13
Vx493 xm493 0 0
Gx493_3 x493 0 u3 0 -7.63577317878425e-08
Rx494 x494 0 1
Fxc494_493 x494 0 Vx493 -139.625080208528
Cx494 x494 xm494 1.4311943973241e-13
Vx494 xm494 0 0
Gx494_3 x494 0 u3 0 1.06614544254188e-05
Rx495 x495 0 1
Fxc495_496 x495 0 Vx496 1165.68249357447
Cx495 x495 xm495 1.49527034425067e-14
Vx495 xm495 0 0
Gx495_3 x495 0 u3 0 -2.63525100931908e-09
Rx496 x496 0 1
Fxc496_495 x496 0 Vx495 -7726.43794539491
Cx496 x496 xm496 1.49527034425067e-14
Vx496 xm496 0 0
Gx496_3 x496 0 u3 0 2.03611033940432e-05
Rx497 x497 0 1
Fxc497_498 x497 0 Vx498 114.595430945885
Cx497 x497 xm497 1.29249231176747e-13
Vx497 xm497 0 0
Gx497_3 x497 0 u3 0 -2.49519938842182e-08
Rx498 x498 0 1
Fxc498_497 x498 0 Vx497 -1091.97923504661
Cx498 x498 xm498 1.29249231176747e-13
Vx498 xm498 0 0
Gx498_3 x498 0 u3 0 2.72470591945763e-05
Rx499 x499 0 1
Fxc499_500 x499 0 Vx500 284.383100144362
Cx499 x499 xm499 2.97577142965506e-14
Vx499 xm499 0 0
Gx499_3 x499 0 u3 0 -1.68205132711153e-09
Rx500 x500 0 1
Fxc500_499 x500 0 Vx499 -8616.76363821543
Cx500 x500 xm500 2.97577142965506e-14
Vx500 xm500 0 0
Gx500_3 x500 0 u3 0 1.44938387130667e-05
Rx501 x501 0 1
Fxc501_502 x501 0 Vx502 58.4925413417388
Cx501 x501 xm501 3.66480875628994e-13
Vx501 xm501 0 0
Gx501_3 x501 0 u3 0 -2.57724827584965e-07
Rx502 x502 0 1
Fxc502_501 x502 0 Vx501 -286.293962175027
Cx502 x502 xm502 3.66480875628994e-13
Vx502 xm502 0 0
Gx502_3 x502 0 u3 0 7.37850620401751e-05
Rx503 x503 0 1
Fxc503_504 x503 0 Vx504 135.422763228254
Cx503 x503 xm503 1.55725403798337e-13
Vx503 xm503 0 0
Gx503_3 x503 0 u3 0 -3.83105520570632e-08
Rx504 x504 0 1
Fxc504_503 x504 0 Vx503 -713.758778224897
Cx504 x504 xm504 1.55725403798336e-13
Vx504 xm504 0 0
Gx504_3 x504 0 u3 0 2.73444928293708e-05
Rx505 x505 0 1
Fxc505_506 x505 0 Vx506 1045.22363096954
Cx505 x505 xm505 2.70690945024366e-14
Vx505 xm505 0 0
Gx505_3 x505 0 u3 0 -4.01925347342828e-09
Rx506 x506 0 1
Fxc506_505 x506 0 Vx505 -3358.34736013361
Cx506 x506 xm506 2.70690945024366e-14
Vx506 xm506 0 0
Gx506_3 x506 0 u3 0 1.34980492921957e-05
Rx507 x507 0 1
Fxc507_508 x507 0 Vx508 350.993797642463
Cx507 x507 xm507 1.05947857159888e-13
Vx507 xm507 0 0
Gx507_3 x507 0 u3 0 -1.31111013672106e-08
Rx508 x508 0 1
Fxc508_507 x508 0 Vx507 -626.451833076192
Cx508 x508 xm508 1.05947857159888e-13
Vx508 xm508 0 0
Gx508_3 x508 0 u3 0 8.21347348513684e-06
Rx509 x509 0 1
Fxc509_510 x509 0 Vx510 160.303007903125
Cx509 x509 xm509 8.05411899100067e-14
Vx509 xm509 0 0
Gx509_3 x509 0 u3 0 -4.21618454311811e-09
Rx510 x510 0 1
Fxc510_509 x510 0 Vx509 -2645.56235269805
Cx510 x510 xm510 8.05411899100067e-14
Vx510 xm510 0 0
Gx510_3 x510 0 u3 0 1.11541790993007e-05
Rx511 x511 0 1
Fxc511_512 x511 0 Vx512 112.273308245124
Cx511 x511 xm511 2.77463484357731e-13
Vx511 xm511 0 0
Gx511_3 x511 0 u3 0 -1.35534247607712e-07
Rx512 x512 0 1
Fxc512_511 x512 0 Vx511 -329.637333614772
Cx512 x512 xm512 2.77463484357731e-13
Vx512 xm512 0 0
Gx512_3 x512 0 u3 0 4.46771479948904e-05
Rx513 x513 0 1
Cx513 x513 0 1.26327330229509e-10
Gx513_3 x513 0 u3 0 -2.59585350182602
Rx514 x514 0 1
Fxc514_515 x514 0 Vx515 252.083208172213
Cx514 x514 xm514 1.99280702854811e-13
Vx514 xm514 0 0
Gx514_3 x514 0 u3 0 -8.04731413788348e-08
Rx515 x515 0 1
Fxc515_514 x515 0 Vx514 -297.932217868013
Cx515 x515 xm515 1.99280702854811e-13
Vx515 xm515 0 0
Gx515_3 x515 0 u3 0 2.39755414898024e-05
Rx516 x516 0 1
Fxc516_517 x516 0 Vx517 1800.42430581648
Cx516 x516 xm516 3.34725367390173e-14
Vx516 xm516 0 0
Gx516_3 x516 0 u3 0 -9.82260423746157e-09
Rx517 x517 0 1
Fxc517_516 x517 0 Vx516 -1560.76028632532
Cx517 x517 xm517 3.34725367390174e-14
Vx517 xm517 0 0
Gx517_3 x517 0 u3 0 1.53307306021209e-05
Rx518 x518 0 1
Fxc518_519 x518 0 Vx519 198.926769517262
Cx518 x518 xm518 1.20981905835219e-12
Vx518 xm518 0 0
Gx518_3 x518 0 u3 0 -9.0989259745268e-06
Rx519 x519 0 1
Fxc519_518 x519 0 Vx518 -11.1735515816997
Cx519 x519 xm519 1.20981905835219e-12
Vx519 xm519 0 0
Gx519_3 x519 0 u3 0 0.000101667318714442
Rx520 x520 0 1
Fxc520_521 x520 0 Vx521 104.874561872073
Cx520 x520 xm520 2.41747187333388e-13
Vx520 xm520 0 0
Gx520_3 x520 0 u3 0 -6.36316459786105e-08
Rx521 x521 0 1
Fxc521_520 x521 0 Vx520 -573.857554438737
Cx521 x521 xm521 2.41747187333388e-13
Vx521 xm521 0 0
Gx521_3 x521 0 u3 0 3.65155007461969e-05
Rx522 x522 0 1
Fxc522_523 x522 0 Vx523 407.101920126474
Cx522 x522 xm522 6.05595987313277e-13
Vx522 xm522 0 0
Gx522_3 x522 0 u3 0 -1.68991851430627e-06
Rx523 x523 0 1
Fxc523_522 x523 0 Vx522 -24.093257535365
Cx523 x523 xm523 6.05595987313277e-13
Vx523 xm523 0 0
Gx523_3 x523 0 u3 0 4.07156419789623e-05
Rx524 x524 0 1
Fxc524_525 x524 0 Vx525 32.0989041139797
Cx524 x524 xm524 4.27273098109608e-12
Vx524 xm524 0 0
Gx524_3 x524 0 u3 0 -0.000328356064243211
Rx525 x525 0 1
Fxc525_524 x525 0 Vx524 -7.17422795018132
Cx525 x525 xm525 4.27273098109608e-12
Vx525 xm525 0 0
Gx525_3 x525 0 u3 0 0.00235570125370518
Rx526 x526 0 1
Fxc526_527 x526 0 Vx527 251.022079360786
Cx526 x526 xm526 2.2113064440014e-13
Vx526 xm526 0 0
Gx526_3 x526 0 u3 0 -4.78052956120523e-08
Rx527 x527 0 1
Fxc527_526 x527 0 Vx526 -318.301722875481
Cx527 x527 xm527 2.2113064440014e-13
Vx527 xm527 0 0
Gx527_3 x527 0 u3 0 1.52165079558879e-05
Rx528 x528 0 1
Fxc528_529 x528 0 Vx529 396.967700227608
Cx528 x528 xm528 3.84635353963742e-13
Vx528 xm528 0 0
Gx528_3 x528 0 u3 0 -3.61360578199969e-07
Rx529 x529 0 1
Fxc529_528 x529 0 Vx528 -69.8872775465159
Cx529 x529 xm529 3.84635353963742e-13
Vx529 xm529 0 0
Gx529_3 x529 0 u3 0 2.52545070230307e-05
Rx530 x530 0 1
Fxc530_531 x530 0 Vx531 22.6809205576968
Cx530 x530 xm530 1.31174697600352e-12
Vx530 xm530 0 0
Gx530_3 x530 0 u3 0 -8.04233689743648e-06
Rx531 x531 0 1
Fxc531_530 x531 0 Vx530 -111.763914440243
Cx531 x531 xm531 1.31174697600352e-12
Vx531 xm531 0 0
Gx531_3 x531 0 u3 0 0.000898843052904699
Rx532 x532 0 1
Fxc532_533 x532 0 Vx533 61.9466514286328
Cx532 x532 xm532 6.73245820833979e-13
Vx532 xm532 0 0
Gx532_3 x532 0 u3 0 -1.42132500176586e-06
Rx533 x533 0 1
Fxc533_532 x533 0 Vx532 -158.080115886001
Cx533 x533 xm533 6.73245820833979e-13
Vx533 xm533 0 0
Gx533_3 x533 0 u3 0 0.000224683220990817
Rx534 x534 0 1
Fxc534_535 x534 0 Vx535 88.761622448351
Cx534 x534 xm534 5.84808784752663e-13
Vx534 xm534 0 0
Gx534_3 x534 0 u3 0 -3.07835781594304e-07
Rx535 x535 0 1
Fxc535_534 x535 0 Vx534 -161.172770138999
Cx535 x535 xm535 5.84808784752663e-13
Vx535 xm535 0 0
Gx535_3 x535 0 u3 0 4.96147456674578e-05
Rx536 x536 0 1
Fxc536_537 x536 0 Vx537 446.895818201252
Cx536 x536 xm536 1.79416446898388e-13
Vx536 xm536 0 0
Gx536_3 x536 0 u3 0 -3.05299701665407e-08
Rx537 x537 0 1
Fxc537_536 x537 0 Vx536 -371.47537960666
Cx537 x537 xm537 1.79416446898388e-13
Vx537 xm537 0 0
Gx537_3 x537 0 u3 0 1.13411322569957e-05
Rx538 x538 0 1
Fxc538_539 x538 0 Vx539 44.7002949791091
Cx538 x538 xm538 9.55321996041439e-13
Vx538 xm538 0 0
Gx538_3 x538 0 u3 0 -8.51921739719417e-07
Rx539 x539 0 1
Fxc539_538 x539 0 Vx538 -143.127440418855
Cx539 x539 xm539 9.55321996041439e-13
Vx539 xm539 0 0
Gx539_3 x539 0 u3 0 0.000121933378043218
Rx540 x540 0 1
Fxc540_541 x540 0 Vx541 40.8618647776235
Cx540 x540 xm540 4.22656817502044e-13
Vx540 xm540 0 0
Gx540_3 x540 0 u3 0 -5.91736740015496e-08
Rx541 x541 0 1
Fxc541_540 x541 0 Vx540 -828.508697954216
Cx541 x541 xm541 4.22656817502044e-13
Vx541 xm541 0 0
Gx541_3 x541 0 u3 0 4.90259036001911e-05
Rx542 x542 0 1
Fxc542_543 x542 0 Vx543 16.666037386787
Cx542 x542 xm542 2.32688864615857e-12
Vx542 xm542 0 0
Gx542_3 x542 0 u3 0 -5.55735447114352e-06
Rx543 x543 0 1
Fxc543_542 x543 0 Vx542 -73.4976540688041
Cx543 x543 xm543 2.32688864615857e-12
Vx543 xm543 0 0
Gx543_3 x543 0 u3 0 0.000408452516457828
Rx544 x544 0 1
Fxc544_545 x544 0 Vx545 275.731015986248
Cx544 x544 xm544 2.24826805546157e-13
Vx544 xm544 0 0
Gx544_3 x544 0 u3 0 -2.44978803822432e-08
Rx545 x545 0 1
Fxc545_544 x545 0 Vx544 -477.948940106319
Cx545 x545 xm545 2.24826805546157e-13
Vx545 xm545 0 0
Gx545_3 x545 0 u3 0 1.17087359635445e-05
Rx546 x546 0 1
Fxc546_547 x546 0 Vx547 170.325190171075
Cx546 x546 xm546 7.62490228495289e-13
Vx546 xm546 0 0
Gx546_3 x546 0 u3 0 -4.68301929755252e-07
Rx547 x547 0 1
Fxc547_546 x547 0 Vx546 -76.1501102886457
Cx547 x547 xm547 7.62490228495289e-13
Vx547 xm547 0 0
Gx547_3 x547 0 u3 0 3.5661243599248e-05
Rx548 x548 0 1
Fxc548_549 x548 0 Vx549 175.491138237085
Cx548 x548 xm548 3.12815339647046e-13
Vx548 xm548 0 0
Gx548_3 x548 0 u3 0 -3.36640336768607e-08
Rx549 x549 0 1
Fxc549_548 x549 0 Vx548 -477.981887976349
Cx549 x549 xm549 3.12815339647046e-13
Vx549 xm549 0 0
Gx549_3 x549 0 u3 0 1.60907983737653e-05
Rx550 x550 0 1
Fxc550_551 x550 0 Vx551 114.866361989283
Cx550 x550 xm550 1.21980473796757e-12
Vx550 xm550 0 0
Gx550_3 x550 0 u3 0 -1.01320363603094e-06
Rx551 x551 0 1
Fxc551_550 x551 0 Vx550 -50.427418100891
Cx551 x551 xm551 1.21980473796757e-12
Vx551 xm551 0 0
Gx551_3 x551 0 u3 0 5.10932433754751e-05
Rx552 x552 0 1
Fxc552_553 x552 0 Vx553 1.39206128507602
Cx552 x552 xm552 6.30927595670662e-12
Vx552 xm552 0 0
Gx552_3 x552 0 u3 0 -8.98083089172031e-06
Rx553 x553 0 1
Fxc553_552 x553 0 Vx552 -183.870533718947
Cx553 x553 xm553 6.30927595670662e-12
Vx553 xm553 0 0
Gx553_3 x553 0 u3 0 0.00165131016930022
Rx554 x554 0 1
Fxc554_555 x554 0 Vx555 7300.5158679474
Cx554 x554 xm554 5.94898906330198e-14
Vx554 xm554 0 0
Gx554_3 x554 0 u3 0 -2.55150886013717e-08
Rx555 x555 0 1
Fxc555_554 x555 0 Vx554 -386.090744907659
Cx555 x555 xm555 5.94898906330198e-14
Vx555 xm555 0 0
Gx555_3 x555 0 u3 0 9.85113956448853e-06
Rx556 x556 0 1
Fxc556_557 x556 0 Vx557 310.423791490136
Cx556 x556 xm556 1.88629779420802e-12
Vx556 xm556 0 0
Gx556_3 x556 0 u3 0 -4.32910166613114e-06
Rx557 x557 0 1
Fxc557_556 x557 0 Vx556 -9.88317802502896
Cx557 x557 xm557 1.88629779420802e-12
Vx557 xm557 0 0
Gx557_3 x557 0 u3 0 4.27852824548235e-05
Rx558 x558 0 1
Fxc558_559 x558 0 Vx559 10.5204245444202
Cx558 x558 xm558 2.53255697284169e-12
Vx558 xm558 0 0
Gx558_3 x558 0 u3 0 -1.64852405200949e-06
Rx559 x559 0 1
Fxc559_558 x559 0 Vx558 -190.3051330805
Cx559 x559 xm559 2.53255697284169e-12
Vx559 xm559 0 0
Gx559_3 x559 0 u3 0 0.000313722589104071
Rx560 x560 0 1
Fxc560_561 x560 0 Vx561 13.3125510454916
Cx560 x560 xm560 1.07068178225324e-12
Vx560 xm560 0 0
Gx560_3 x560 0 u3 0 -1.07540721902096e-07
Rx561 x561 0 1
Fxc561_560 x561 0 Vx560 -899.540343605639
Cx561 x561 xm561 1.07068178225324e-12
Vx561 xm561 0 0
Gx561_3 x561 0 u3 0 9.673721793141e-05
Rx562 x562 0 1
Cx562 x562 0 5.22190407222509e-10
Gx562_3 x562 0 u3 0 -0.290427634715475
Rx563 x563 0 1
Fxc563_564 x563 0 Vx564 85.5040310330202
Cx563 x563 xm563 1.10121754249303e-12
Vx563 xm563 0 0
Gx563_3 x563 0 u3 0 -2.89192738066707e-07
Rx564 x564 0 1
Fxc564_563 x564 0 Vx563 -161.253515946278
Cx564 x564 xm564 1.10121754249303e-12
Vx564 xm564 0 0
Gx564_3 x564 0 u3 0 4.66333457993875e-05
Rx565 x565 0 1
Fxc565_566 x565 0 Vx566 176.511581021896
Cx565 x565 xm565 1.35840059784609e-12
Vx565 xm565 0 0
Gx565_3 x565 0 u3 0 -5.32906731466139e-07
Rx566 x566 0 1
Fxc566_565 x566 0 Vx565 -58.6605867806999
Cx566 x566 xm566 1.3584005978461e-12
Vx566 xm566 0 0
Gx566_3 x566 0 u3 0 3.12606215671886e-05
Rx567 x567 0 1
Fxc567_568 x567 0 Vx568 7.98835078316539
Cx567 x567 xm567 1.37582820475616e-11
Vx567 xm567 0 0
Gx567_3 x567 0 u3 0 -9.77278180239205e-05
Rx568 x568 0 1
Fxc568_567 x568 0 Vx567 -17.4576478721131
Cx568 x568 xm568 1.37582820475616e-11
Vx568 xm568 0 0
Gx568_3 x568 0 u3 0 0.00170609783437155
Rx569 x569 0 1
Fxc569_570 x569 0 Vx570 18.8506926539648
Cx569 x569 xm569 2.55525080407755e-12
Vx569 xm569 0 0
Gx569_3 x569 0 u3 0 -2.11860908543465e-06
Rx570 x570 0 1
Fxc570_569 x570 0 Vx569 -118.390709457023
Cx570 x570 xm570 2.55525080407755e-12
Vx570 xm570 0 0
Gx570_3 x570 0 u3 0 0.000250823632686703
Rx571 x571 0 1
Fxc571_572 x571 0 Vx572 17.5741111749443
Cx571 x571 xm571 3.52048110577458e-12
Vx571 xm571 0 0
Gx571_3 x571 0 u3 0 -2.20224038937497e-06
Rx572 x572 0 1
Fxc572_571 x572 0 Vx571 -100.451259503632
Cx572 x572 xm572 3.52048110577458e-12
Vx572 xm572 0 0
Gx572_3 x572 0 u3 0 0.000221217820842485
Rx573 x573 0 1
Fxc573_574 x573 0 Vx574 1.67555439705407
Cx573 x573 xm573 8.01925764208566e-11
Vx573 xm573 0 0
Gx573_3 x573 0 u3 0 -0.00778236392221692
Rx574 x574 0 1
Fxc574_573 x574 0 Vx573 -4.66181176204352
Cx574 x574 xm574 8.01925764208566e-11
Vx574 xm574 0 0
Gx574_3 x574 0 u3 0 0.036279915669094
Rx575 x575 0 1
Fxc575_576 x575 0 Vx576 17.4505717652724
Cx575 x575 xm575 1.34818539204243e-12
Vx575 xm575 0 0
Gx575_3 x575 0 u3 0 -5.90853364881975e-08
Rx576 x576 0 1
Fxc576_575 x576 0 Vx575 -864.835545863289
Cx576 x576 xm576 1.34818539204243e-12
Vx576 xm576 0 0
Gx576_3 x576 0 u3 0 5.10990992342864e-05
Rx577 x577 0 1
Fxc577_578 x577 0 Vx578 2.33462606056593
Cx577 x577 xm577 2.60286578934868e-10
Vx577 xm577 0 0
Gx577_3 x577 0 u3 0 -0.0311857849870516
Rx578 x578 0 1
Fxc578_577 x578 0 Vx577 -1.26083198071759
Cx578 x578 xm578 2.60286578934868e-10
Vx578 xm578 0 0
Gx578_3 x578 0 u3 0 0.039320035055457
Rx579 x579 0 1
Fxc579_580 x579 0 Vx580 25.5625489869627
Cx579 x579 xm579 1.94992797826926e-12
Vx579 xm579 0 0
Gx579_3 x579 0 u3 0 -1.85522653561035e-07
Rx580 x580 0 1
Fxc580_579 x580 0 Vx579 -352.247523794223
Cx580 x580 xm580 1.94992797826926e-12
Vx580 xm580 0 0
Gx580_3 x580 0 u3 0 6.53498953246079e-05
Rx581 x581 0 1
Fxc581_582 x581 0 Vx582 129.58703747971
Cx581 x581 xm581 2.33413529363335e-12
Vx581 xm581 0 0
Gx581_3 x581 0 u3 0 -2.32279426491235e-07
Rx582 x582 0 1
Fxc582_581 x582 0 Vx581 -125.985228933684
Cx582 x582 xm582 2.33413529363335e-12
Vx582 xm582 0 0
Gx582_3 x582 0 u3 0 2.9263776723083e-05
Rx583 x583 0 1
Fxc583_584 x583 0 Vx584 6.15575630366068
Cx583 x583 xm583 1.72271737747677e-11
Vx583 xm583 0 0
Gx583_3 x583 0 u3 0 -3.0045611333238e-05
Rx584 x584 0 1
Fxc584_583 x584 0 Vx583 -33.8490622197189
Cx584 x584 xm584 1.72271737747677e-11
Vx584 xm584 0 0
Gx584_3 x584 0 u3 0 0.00101701576744826
Rx585 x585 0 1
Fxc585_586 x585 0 Vx586 315.313297299494
Cx585 x585 xm585 3.38373728470339e-12
Vx585 xm585 0 0
Gx585_3 x585 0 u3 0 -1.84085111398413e-06
Rx586 x586 0 1
Fxc586_585 x586 0 Vx585 -11.805776931499
Cx586 x586 xm586 3.38373728470339e-12
Vx586 xm586 0 0
Gx586_3 x586 0 u3 0 2.17326776157981e-05
Rx587 x587 0 1
Fxc587_588 x587 0 Vx588 73.8109027147112
Cx587 x587 xm587 5.83456226648167e-12
Vx587 xm587 0 0
Gx587_3 x587 0 u3 0 -9.8188727258034e-07
Rx588 x588 0 1
Fxc588_587 x588 0 Vx587 -57.845737290184
Cx588 x588 xm588 5.83456226648167e-12
Vx588 xm588 0 0
Gx588_3 x588 0 u3 0 5.67979932182577e-05
Rx589 x589 0 1
Fxc589_590 x589 0 Vx590 16.7935180797451
Cx589 x589 xm589 3.71913677806581e-11
Vx589 xm589 0 0
Gx589_3 x589 0 u3 0 -0.000870584594886927
Rx590 x590 0 1
Fxc590_589 x590 0 Vx589 -11.2719975033048
Cx590 x590 xm590 3.71913677806581e-11
Vx590 xm590 0 0
Gx590_3 x590 0 u3 0 0.00981322737998107
Rx591 x591 0 1
Fxc591_592 x591 0 Vx592 15.4860101676856
Cx591 x591 xm591 3.43647746350443e-11
Vx591 xm591 0 0
Gx591_3 x591 0 u3 0 -0.000659309033592774
Rx592 x592 0 1
Fxc592_591 x592 0 Vx591 -14.2465477032417
Cx592 x592 xm592 3.43647746350443e-11
Vx592 xm592 0 0
Gx592_3 x592 0 u3 0 0.00939287759825765
Rx593 x593 0 1
Fxc593_594 x593 0 Vx594 6.85757771599204
Cx593 x593 xm593 1.92407202503742e-10
Vx593 xm593 0 0
Gx593_3 x593 0 u3 0 -0.000480239816844695
Rx594 x594 0 1
Fxc594_593 x594 0 Vx593 -3.57511563582002
Cx594 x594 xm594 1.92407202503742e-10
Vx594 xm594 0 0
Gx594_3 x594 0 u3 0 0.00171691287814481
Rx595 x595 0 1
Fxc595_596 x595 0 Vx596 797.185649131755
Cx595 x595 xm595 8.89563374249556e-13
Vx595 xm595 0 0
Gx595_3 x595 0 u3 0 -1.64347868555196e-07
Rx596 x596 0 1
Fxc596_595 x596 0 Vx595 -93.5216567317908
Cx596 x596 xm596 8.89563374249556e-13
Vx596 xm596 0 0
Gx596_3 x596 0 u3 0 1.53700849476205e-05
Rx597 x597 0 1
Fxc597_598 x597 0 Vx598 1.00445350908454
Cx597 x597 xm597 1.38719414317867e-09
Vx597 xm597 0 0
Gx597_3 x597 0 u3 0 -0.0295648309716011
Rx598 x598 0 1
Fxc598_597 x598 0 Vx597 -0.579938038060297
Cx598 x598 xm598 1.38719414317867e-09
Vx598 xm598 0 0
Gx598_3 x598 0 u3 0 0.0171457700692546
Rx599 x599 0 1
Cx599 x599 0 4.58826427740312e-07
Gx599_3 x599 0 u3 0 -0.585742874013833
Rx600 x600 0 1
Cx600 x600 0 7.53723517430562e-08
Gx600_3 x600 0 u3 0 -0.291148167471246
Gyc1_1 y1 0 x1 0 -1
Gyc1_2 y1 0 x2 0 1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 1
Gyc1_5 y1 0 x5 0 -0.825114395183513
Gyc1_6 y1 0 x6 0 1
Gyc1_7 y1 0 x7 0 -1
Gyc1_8 y1 0 x8 0 1
Gyc1_9 y1 0 x9 0 -1
Gyc1_10 y1 0 x10 0 -1
Gyc1_11 y1 0 x11 0 -1
Gyc1_12 y1 0 x12 0 0.109193707790164
Gyc1_13 y1 0 x13 0 -1
Gyc1_14 y1 0 x14 0 -1
Gyc1_15 y1 0 x15 0 1
Gyc1_16 y1 0 x16 0 -1
Gyc1_17 y1 0 x17 0 1
Gyc1_18 y1 0 x18 0 -1
Gyc1_19 y1 0 x19 0 1
Gyc1_20 y1 0 x20 0 1
Gyc1_21 y1 0 x21 0 1
Gyc1_22 y1 0 x22 0 1
Gyc1_23 y1 0 x23 0 -1
Gyc1_24 y1 0 x24 0 1
Gyc1_25 y1 0 x25 0 -1
Gyc1_26 y1 0 x26 0 1
Gyc1_27 y1 0 x27 0 1
Gyc1_28 y1 0 x28 0 -1
Gyc1_29 y1 0 x29 0 -1
Gyc1_30 y1 0 x30 0 1
Gyc1_31 y1 0 x31 0 -1
Gyc1_32 y1 0 x32 0 -1
Gyc1_33 y1 0 x33 0 1
Gyc1_34 y1 0 x34 0 1
Gyc1_35 y1 0 x35 0 1
Gyc1_36 y1 0 x36 0 -1
Gyc1_37 y1 0 x37 0 -1
Gyc1_38 y1 0 x38 0 1
Gyc1_39 y1 0 x39 0 1
Gyc1_40 y1 0 x40 0 -1
Gyc1_41 y1 0 x41 0 1
Gyc1_42 y1 0 x42 0 -1
Gyc1_43 y1 0 x43 0 0.684147443107
Gyc1_44 y1 0 x44 0 1
Gyc1_45 y1 0 x45 0 1
Gyc1_46 y1 0 x46 0 1
Gyc1_47 y1 0 x47 0 1
Gyc1_48 y1 0 x48 0 1
Gyc1_49 y1 0 x49 0 1
Gyc1_50 y1 0 x50 0 1
Gyc1_51 y1 0 x51 0 -1
Gyc1_52 y1 0 x52 0 1
Gyc1_53 y1 0 x53 0 -1
Gyc1_54 y1 0 x54 0 -1
Gyc1_55 y1 0 x55 0 -1
Gyc1_56 y1 0 x56 0 1
Gyc1_57 y1 0 x57 0 -1
Gyc1_58 y1 0 x58 0 -1
Gyc1_59 y1 0 x59 0 -1
Gyc1_60 y1 0 x60 0 -1
Gyc1_61 y1 0 x61 0 1
Gyc1_62 y1 0 x62 0 -0.508197051165551
Gyc1_63 y1 0 x63 0 -1
Gyc1_64 y1 0 x64 0 -1
Gyc1_65 y1 0 x65 0 0.355570912418791
Gyc1_66 y1 0 x66 0 1
Gyc1_67 y1 0 x67 0 1
Gyc1_68 y1 0 x68 0 1
Gyc1_69 y1 0 x69 0 -1
Gyc1_70 y1 0 x70 0 1
Gyc1_71 y1 0 x71 0 -1
Gyc1_72 y1 0 x72 0 0.981851444758819
Gyc1_73 y1 0 x73 0 -1
Gyc1_74 y1 0 x74 0 -1
Gyc1_75 y1 0 x75 0 -1
Gyc1_76 y1 0 x76 0 -1
Gyc1_77 y1 0 x77 0 1
Gyc1_78 y1 0 x78 0 -1
Gyc1_79 y1 0 x79 0 -1
Gyc1_80 y1 0 x80 0 -1
Gyc1_81 y1 0 x81 0 -1
Gyc1_82 y1 0 x82 0 1
Gyc1_83 y1 0 x83 0 -1
Gyc1_84 y1 0 x84 0 0.37928566566302
Gyc1_85 y1 0 x85 0 0.970032171227361
Gyc1_86 y1 0 x86 0 -1
Gyc1_87 y1 0 x87 0 1
Gyc1_88 y1 0 x88 0 -1
Gyc1_89 y1 0 x89 0 1
Gyc1_90 y1 0 x90 0 -1
Gyc1_91 y1 0 x91 0 1
Gyc1_92 y1 0 x92 0 -1
Gyc1_93 y1 0 x93 0 1
Gyc1_94 y1 0 x94 0 1
Gyc1_95 y1 0 x95 0 -1
Gyc1_96 y1 0 x96 0 1
Gyc1_97 y1 0 x97 0 0.305778402553825
Gyc1_98 y1 0 x98 0 1
Gyc1_99 y1 0 x99 0 -1
Gyc1_100 y1 0 x100 0 1
Gyc1_101 y1 0 x101 0 -1
Gyc1_102 y1 0 x102 0 1
Gyc1_103 y1 0 x103 0 -1
Gyc1_104 y1 0 x104 0 0.819980794754496
Gyc1_105 y1 0 x105 0 1
Gyc1_106 y1 0 x106 0 -1
Gyc1_107 y1 0 x107 0 -1
Gyc1_108 y1 0 x108 0 -1
Gyc1_109 y1 0 x109 0 1
Gyc1_110 y1 0 x110 0 -1
Gyc1_111 y1 0 x111 0 1
Gyc1_112 y1 0 x112 0 -1
Gyc1_113 y1 0 x113 0 1
Gyc1_114 y1 0 x114 0 1
Gyc1_115 y1 0 x115 0 1
Gyc1_116 y1 0 x116 0 1
Gyc1_117 y1 0 x117 0 1
Gyc1_118 y1 0 x118 0 1
Gyc1_119 y1 0 x119 0 1
Gyc1_120 y1 0 x120 0 -1
Gyc1_121 y1 0 x121 0 1
Gyc1_122 y1 0 x122 0 1
Gyc1_123 y1 0 x123 0 1
Gyc1_124 y1 0 x124 0 1
Gyc1_125 y1 0 x125 0 1
Gyc1_126 y1 0 x126 0 -1
Gyc1_127 y1 0 x127 0 1
Gyc1_128 y1 0 x128 0 -1
Gyc1_129 y1 0 x129 0 -1
Gyc1_130 y1 0 x130 0 1
Gyc1_131 y1 0 x131 0 -1
Gyc1_132 y1 0 x132 0 -1
Gyc1_133 y1 0 x133 0 1
Gyc1_134 y1 0 x134 0 1
Gyc1_135 y1 0 x135 0 -1
Gyc1_136 y1 0 x136 0 1
Gyc1_137 y1 0 x137 0 1
Gyc1_138 y1 0 x138 0 -1
Gyc1_139 y1 0 x139 0 1
Gyc1_140 y1 0 x140 0 -1
Gyc1_141 y1 0 x141 0 1
Gyc1_142 y1 0 x142 0 -1
Gyc1_143 y1 0 x143 0 1
Gyc1_144 y1 0 x144 0 1
Gyc1_145 y1 0 x145 0 -1
Gyc1_146 y1 0 x146 0 -1
Gyc1_147 y1 0 x147 0 -1
Gyc1_148 y1 0 x148 0 -1
Gyc1_149 y1 0 x149 0 -1
Gyc1_150 y1 0 x150 0 -1
Gyc1_151 y1 0 x151 0 -1
Gyc1_152 y1 0 x152 0 1
Gyc1_153 y1 0 x153 0 -1
Gyc1_154 y1 0 x154 0 -1
Gyc1_155 y1 0 x155 0 1
Gyc1_156 y1 0 x156 0 -1
Gyc1_157 y1 0 x157 0 -1
Gyc1_158 y1 0 x158 0 1
Gyc1_159 y1 0 x159 0 -1
Gyc1_160 y1 0 x160 0 1
Gyc1_161 y1 0 x161 0 -1
Gyc1_162 y1 0 x162 0 -1
Gyc1_163 y1 0 x163 0 1
Gyc1_164 y1 0 x164 0 -1
Gyc1_165 y1 0 x165 0 1
Gyc1_166 y1 0 x166 0 1
Gyc1_167 y1 0 x167 0 1
Gyc1_168 y1 0 x168 0 1
Gyc1_169 y1 0 x169 0 -1
Gyc1_170 y1 0 x170 0 -1
Gyc1_171 y1 0 x171 0 1
Gyc1_172 y1 0 x172 0 1
Gyc1_173 y1 0 x173 0 -1
Gyc1_174 y1 0 x174 0 1
Gyc1_175 y1 0 x175 0 1
Gyc1_176 y1 0 x176 0 -1
Gyc1_177 y1 0 x177 0 -1
Gyc1_178 y1 0 x178 0 -1
Gyc1_179 y1 0 x179 0 -1
Gyc1_180 y1 0 x180 0 1
Gyc1_181 y1 0 x181 0 1
Gyc1_182 y1 0 x182 0 1
Gyc1_183 y1 0 x183 0 1
Gyc1_184 y1 0 x184 0 -1
Gyc1_185 y1 0 x185 0 -1
Gyc1_186 y1 0 x186 0 -1
Gyc1_187 y1 0 x187 0 -1
Gyc1_188 y1 0 x188 0 -1
Gyc1_189 y1 0 x189 0 1
Gyc1_190 y1 0 x190 0 -1
Gyc1_191 y1 0 x191 0 -1
Gyc1_192 y1 0 x192 0 1
Gyc1_193 y1 0 x193 0 -1
Gyc1_194 y1 0 x194 0 -1
Gyc1_195 y1 0 x195 0 1
Gyc1_196 y1 0 x196 0 1
Gyc1_197 y1 0 x197 0 1
Gyc1_198 y1 0 x198 0 -1
Gyc1_199 y1 0 x199 0 1
Gyc1_200 y1 0 x200 0 1
Gyc1_201 y1 0 x201 0 -0.299981825501131
Gyc1_202 y1 0 x202 0 -0.338380278115099
Gyc1_203 y1 0 x203 0 0.161234663785178
Gyc1_204 y1 0 x204 0 -0.416754089085469
Gyc1_205 y1 0 x205 0 -0.211597147135213
Gyc1_206 y1 0 x206 0 0.0673680577069801
Gyc1_207 y1 0 x207 0 -0.239095187988776
Gyc1_208 y1 0 x208 0 -0.0806496060198992
Gyc1_209 y1 0 x209 0 2.08176977078619e-05
Gyc1_210 y1 0 x210 0 0.336218635416246
Gyc1_211 y1 0 x211 0 0.0250700361537084
Gyc1_212 y1 0 x212 0 -0.325758981693414
Gyc1_213 y1 0 x213 0 0.245638738610268
Gyc1_214 y1 0 x214 0 -0.359511426689917
Gyc1_215 y1 0 x215 0 -0.296369809668037
Gyc1_216 y1 0 x216 0 0.437260047218514
Gyc1_217 y1 0 x217 0 0.527871568902346
Gyc1_218 y1 0 x218 0 -0.177091830392313
Gyc1_219 y1 0 x219 0 0.192708785181276
Gyc1_220 y1 0 x220 0 -0.0672343614661195
Gyc1_221 y1 0 x221 0 -0.161262169254523
Gyc1_222 y1 0 x222 0 0.0972509552719221
Gyc1_223 y1 0 x223 0 0.18555891948954
Gyc1_224 y1 0 x224 0 0.0563857347534709
Gyc1_225 y1 0 x225 0 0.11496965583329
Gyc1_226 y1 0 x226 0 -0.418551442632015
Gyc1_227 y1 0 x227 0 -1
Gyc1_228 y1 0 x228 0 0.0597051321983344
Gyc1_229 y1 0 x229 0 -0.335291817258667
Gyc1_230 y1 0 x230 0 -1
Gyc1_231 y1 0 x231 0 0.309700466712937
Gyc1_232 y1 0 x232 0 -0.491229223138836
Gyc1_233 y1 0 x233 0 0.289238995506214
Gyc1_234 y1 0 x234 0 -0.210090124077598
Gyc1_235 y1 0 x235 0 0.0521867867329834
Gyc1_236 y1 0 x236 0 0.0825645763741608
Gyc1_237 y1 0 x237 0 -1
Gyc1_238 y1 0 x238 0 -0.0893370889871398
Gyc1_239 y1 0 x239 0 -0.517440397586779
Gyc1_240 y1 0 x240 0 -0.378601858739769
Gyc1_241 y1 0 x241 0 -1
Gyc1_242 y1 0 x242 0 1
Gyc1_243 y1 0 x243 0 -1
Gyc1_244 y1 0 x244 0 0.749467535986598
Gyc1_245 y1 0 x245 0 0.106482311790286
Gyc1_246 y1 0 x246 0 -0.127183877937944
Gyc1_247 y1 0 x247 0 -1
Gyc1_248 y1 0 x248 0 -0.179105118986054
Gyc1_249 y1 0 x249 0 -0.270774014250882
Gyc1_250 y1 0 x250 0 0.179844332358671
Gyc1_251 y1 0 x251 0 -0.113470703707672
Gyc1_252 y1 0 x252 0 0.564909133492989
Gyc1_253 y1 0 x253 0 0.202276157520173
Gyc1_254 y1 0 x254 0 1
Gyc1_255 y1 0 x255 0 -0.248125796719312
Gyc1_256 y1 0 x256 0 -0.223624528449511
Gyc1_257 y1 0 x257 0 1
Gyc1_258 y1 0 x258 0 0.893775507450794
Gyc1_259 y1 0 x259 0 -0.533580315276294
Gyc1_260 y1 0 x260 0 -0.550598301739976
Gyc1_261 y1 0 x261 0 -1
Gyc1_262 y1 0 x262 0 0.372230786352272
Gyc1_263 y1 0 x263 0 0.286042479860404
Gyc1_264 y1 0 x264 0 0.0306461810483885
Gyc1_265 y1 0 x265 0 -1
Gyc1_266 y1 0 x266 0 0.513850327518182
Gyc1_267 y1 0 x267 0 -0.0104507466383546
Gyc1_268 y1 0 x268 0 -1
Gyc1_269 y1 0 x269 0 0.226873353623264
Gyc1_270 y1 0 x270 0 0.00495576456937673
Gyc1_271 y1 0 x271 0 -0.957083887041806
Gyc1_272 y1 0 x272 0 -0.913650505097616
Gyc1_273 y1 0 x273 0 -0.945812253611419
Gyc1_274 y1 0 x274 0 0.16834473949534
Gyc1_275 y1 0 x275 0 1
Gyc1_276 y1 0 x276 0 -0.455510144939363
Gyc1_277 y1 0 x277 0 -0.532672726393711
Gyc1_278 y1 0 x278 0 -0.994963278485022
Gyc1_279 y1 0 x279 0 -0.227403502521678
Gyc1_280 y1 0 x280 0 0.487769927147804
Gyc1_281 y1 0 x281 0 -1
Gyc1_282 y1 0 x282 0 -0.176575330810881
Gyc1_283 y1 0 x283 0 -0.690353149803887
Gyc1_284 y1 0 x284 0 0.945910990538579
Gyc1_285 y1 0 x285 0 0.67342119597286
Gyc1_286 y1 0 x286 0 1
Gyc1_287 y1 0 x287 0 -1
Gyc1_288 y1 0 x288 0 -1
Gyc1_289 y1 0 x289 0 -0.530895256096341
Gyc1_290 y1 0 x290 0 0.410985079249119
Gyc1_291 y1 0 x291 0 0.0376421122795325
Gyc1_292 y1 0 x292 0 -0.275125391665439
Gyc1_293 y1 0 x293 0 -0.813094917956758
Gyc1_294 y1 0 x294 0 -1
Gyc1_295 y1 0 x295 0 -0.158182945036477
Gyc1_296 y1 0 x296 0 0.119082796569836
Gyc1_297 y1 0 x297 0 1
Gyc1_298 y1 0 x298 0 -1
Gyc1_299 y1 0 x299 0 -0.909678762195151
Gyc1_300 y1 0 x300 0 0.0877479946962593
Gyc1_301 y1 0 x301 0 0.598589281830503
Gyc1_302 y1 0 x302 0 -1
Gyc1_303 y1 0 x303 0 -0.56585617793207
Gyc1_304 y1 0 x304 0 -1
Gyc1_305 y1 0 x305 0 0.202046557892802
Gyc1_306 y1 0 x306 0 0.0121479419807996
Gyc1_307 y1 0 x307 0 -0.28865603171026
Gyc1_308 y1 0 x308 0 0.420447025141069
Gyc1_309 y1 0 x309 0 0.761403759158718
Gyc1_310 y1 0 x310 0 -0.272468931870497
Gyc1_311 y1 0 x311 0 -0.345144148428477
Gyc1_312 y1 0 x312 0 1
Gyc1_313 y1 0 x313 0 0.159633118669028
Gyc1_314 y1 0 x314 0 0.834463577878566
Gyc1_315 y1 0 x315 0 0.00832053159830302
Gyc1_316 y1 0 x316 0 -0.146377913233858
Gyc1_317 y1 0 x317 0 -0.075991692065023
Gyc1_318 y1 0 x318 0 0.0391372189273834
Gyc1_319 y1 0 x319 0 0.0311993305858794
Gyc1_320 y1 0 x320 0 0.562329410493961
Gyc1_321 y1 0 x321 0 -0.354198375078342
Gyc1_322 y1 0 x322 0 -0.0938243418868679
Gyc1_323 y1 0 x323 0 -0.0392713643471314
Gyc1_324 y1 0 x324 0 0.138894684549954
Gyc1_325 y1 0 x325 0 -0.0839268331080003
Gyc1_326 y1 0 x326 0 0.482106662615311
Gyc1_327 y1 0 x327 0 1
Gyc1_328 y1 0 x328 0 -0.356801688835079
Gyc1_329 y1 0 x329 0 -0.321488912938395
Gyc1_330 y1 0 x330 0 -0.11896897420225
Gyc1_331 y1 0 x331 0 0.0277313167722724
Gyc1_332 y1 0 x332 0 -0.144367117980879
Gyc1_333 y1 0 x333 0 0.0159546763308784
Gyc1_334 y1 0 x334 0 -0.300523267610652
Gyc1_335 y1 0 x335 0 0.0491586051349686
Gyc1_336 y1 0 x336 0 -0.523769017820648
Gyc1_337 y1 0 x337 0 0.168124817056209
Gyc1_338 y1 0 x338 0 0.147675023555711
Gyc1_339 y1 0 x339 0 0.0238010772046884
Gyc1_340 y1 0 x340 0 -0.3923638938397
Gyc1_341 y1 0 x341 0 -0.184503248031562
Gyc1_342 y1 0 x342 0 -0.0411637628223283
Gyc1_343 y1 0 x343 0 0.0473484481680502
Gyc1_344 y1 0 x344 0 -0.23888928892964
Gyc1_345 y1 0 x345 0 1
Gyc1_346 y1 0 x346 0 -0.337870215719539
Gyc1_347 y1 0 x347 0 0.131048505173842
Gyc1_348 y1 0 x348 0 0.495495370637508
Gyc1_349 y1 0 x349 0 0.250044734583303
Gyc1_350 y1 0 x350 0 -1
Gyc1_351 y1 0 x351 0 0.00399473876892962
Gyc1_352 y1 0 x352 0 -0.723953889890171
Gyc1_353 y1 0 x353 0 0.222584869561298
Gyc1_354 y1 0 x354 0 -0.0369101809668661
Gyc1_355 y1 0 x355 0 -0.177659371635734
Gyc1_356 y1 0 x356 0 0.537837117559654
Gyc1_357 y1 0 x357 0 0.9129358084293
Gyc1_358 y1 0 x358 0 -0.0367447486333831
Gyc1_359 y1 0 x359 0 0.657223673096696
Gyc1_360 y1 0 x360 0 -0.0313186412430128
Gyc1_361 y1 0 x361 0 0.228705311887276
Gyc1_362 y1 0 x362 0 0.000625032963633872
Gyc1_363 y1 0 x363 0 0.371942698663149
Gyc1_364 y1 0 x364 0 -0.185965290754105
Gyc1_365 y1 0 x365 0 -1
Gyc1_366 y1 0 x366 0 -0.0625632661870589
Gyc1_367 y1 0 x367 0 -0.358284106985655
Gyc1_368 y1 0 x368 0 -0.206290930910644
Gyc1_369 y1 0 x369 0 1
Gyc1_370 y1 0 x370 0 0.326491101088017
Gyc1_371 y1 0 x371 0 0.0945379669140505
Gyc1_372 y1 0 x372 0 0.164688427731393
Gyc1_373 y1 0 x373 0 0.0236860500605636
Gyc1_374 y1 0 x374 0 -0.31535533696925
Gyc1_375 y1 0 x375 0 0.266846516148672
Gyc1_376 y1 0 x376 0 0.634990061037226
Gyc1_377 y1 0 x377 0 0.327822861544215
Gyc1_378 y1 0 x378 0 -0.0783964869121525
Gyc1_379 y1 0 x379 0 1
Gyc1_380 y1 0 x380 0 0.00517547235269526
Gyc1_381 y1 0 x381 0 0.321548880220443
Gyc1_382 y1 0 x382 0 -0.0341144152645055
Gyc1_383 y1 0 x383 0 0.107237055336929
Gyc1_384 y1 0 x384 0 0.482383964378154
Gyc1_385 y1 0 x385 0 0.56123527749243
Gyc1_386 y1 0 x386 0 -0.255251535600084
Gyc1_387 y1 0 x387 0 0.761842641545933
Gyc1_388 y1 0 x388 0 0.15599558724823
Gyc1_389 y1 0 x389 0 0.0239083884776266
Gyc1_390 y1 0 x390 0 1
Gyc1_391 y1 0 x391 0 -0.037729937792865
Gyc1_392 y1 0 x392 0 -1
Gyc1_393 y1 0 x393 0 0.949873070727895
Gyc1_394 y1 0 x394 0 0.106039529329614
Gyc1_395 y1 0 x395 0 -0.00797885155341218
Gyc1_396 y1 0 x396 0 -0.0128885710229404
Gyc1_397 y1 0 x397 0 0.210937646262333
Gyc1_398 y1 0 x398 0 1
Gyc1_399 y1 0 x399 0 0.547444894494108
Gyc1_400 y1 0 x400 0 0.249030823190402
Gyc1_401 y1 0 x401 0 -0.136664909944813
Gyc1_402 y1 0 x402 0 0.0873810230941248
Gyc1_403 y1 0 x403 0 0.00346370076459404
Gyc1_404 y1 0 x404 0 0.149587233039287
Gyc1_405 y1 0 x405 0 -0.0755166207833754
Gyc1_406 y1 0 x406 0 0.0567675112501105
Gyc1_407 y1 0 x407 0 -0.355684041495528
Gyc1_408 y1 0 x408 0 -0.0343761826963935
Gyc1_409 y1 0 x409 0 0.0412734703135076
Gyc1_410 y1 0 x410 0 0.0343888179532601
Gyc1_411 y1 0 x411 0 0.0312311883717707
Gyc1_412 y1 0 x412 0 -0.103260192992991
Gyc1_413 y1 0 x413 0 0.0600523572162167
Gyc1_414 y1 0 x414 0 -0.353722212928956
Gyc1_415 y1 0 x415 0 0.264934258693749
Gyc1_416 y1 0 x416 0 -0.203726475435171
Gyc1_417 y1 0 x417 0 0.414787924266247
Gyc1_418 y1 0 x418 0 -0.0686134714752985
Gyc1_419 y1 0 x419 0 0.115561452266108
Gyc1_420 y1 0 x420 0 -0.0251526487558031
Gyc1_421 y1 0 x421 0 -0.0513998753937611
Gyc1_422 y1 0 x422 0 -0.0236922780914371
Gyc1_423 y1 0 x423 0 0.0571323423632484
Gyc1_424 y1 0 x424 0 0.117049135299403
Gyc1_425 y1 0 x425 0 0.116116589159253
Gyc1_426 y1 0 x426 0 0.0838255294158483
Gyc1_427 y1 0 x427 0 0.025705840000176
Gyc1_428 y1 0 x428 0 -0.146101710294838
Gyc1_429 y1 0 x429 0 0.416464302570449
Gyc1_430 y1 0 x430 0 0.0791793734497744
Gyc1_431 y1 0 x431 0 -0.00468220033601162
Gyc1_432 y1 0 x432 0 0.231353168296187
Gyc1_433 y1 0 x433 0 0.00575832525353768
Gyc1_434 y1 0 x434 0 0.136499017315217
Gyc1_435 y1 0 x435 0 0.0106700860758177
Gyc1_436 y1 0 x436 0 -0.0374547238344802
Gyc1_437 y1 0 x437 0 0.0962028184180469
Gyc1_438 y1 0 x438 0 0.0306239441655193
Gyc1_439 y1 0 x439 0 0.179504687230513
Gyc1_440 y1 0 x440 0 0.0406929539890873
Gyc1_441 y1 0 x441 0 0.343082678742437
Gyc1_442 y1 0 x442 0 0.0331784040660736
Gyc1_443 y1 0 x443 0 0.195134446673491
Gyc1_444 y1 0 x444 0 0.167030926078474
Gyc1_445 y1 0 x445 0 -0.0298249905746448
Gyc1_446 y1 0 x446 0 -0.000974075580680787
Gyc1_447 y1 0 x447 0 0.0635824002704673
Gyc1_448 y1 0 x448 0 0.335416389978491
Gyc1_449 y1 0 x449 0 0.0876971539160215
Gyc1_450 y1 0 x450 0 0.00200856611066929
Gyc1_451 y1 0 x451 0 1
Gyc1_452 y1 0 x452 0 0.00580578278600666
Gyc1_453 y1 0 x453 0 0.215045719556532
Gyc1_454 y1 0 x454 0 -0.450225983793795
Gyc1_455 y1 0 x455 0 -0.581371748244701
Gyc1_456 y1 0 x456 0 0.0421403370421942
Gyc1_457 y1 0 x457 0 0.0937468829787875
Gyc1_458 y1 0 x458 0 -0.193968738907952
Gyc1_459 y1 0 x459 0 -0.733980664798448
Gyc1_460 y1 0 x460 0 0.381693545456659
Gyc1_461 y1 0 x461 0 -0.0476111578806983
Gyc1_462 y1 0 x462 0 0.486754771257776
Gyc1_463 y1 0 x463 0 -0.0801811436676284
Gyc1_464 y1 0 x464 0 -0.107502921649585
Gyc1_465 y1 0 x465 0 -0.0661893282981747
Gyc1_466 y1 0 x466 0 0.967719506242129
Gyc1_467 y1 0 x467 0 -0.0398167971042757
Gyc1_468 y1 0 x468 0 -0.282057057441158
Gyc1_469 y1 0 x469 0 -0.213349984789514
Gyc1_470 y1 0 x470 0 0.0332466526023264
Gyc1_471 y1 0 x471 0 -1
Gyc1_472 y1 0 x472 0 0.015610025190561
Gyc1_473 y1 0 x473 0 -0.403248108664061
Gyc1_474 y1 0 x474 0 1
Gyc1_475 y1 0 x475 0 0.212862514215524
Gyc1_476 y1 0 x476 0 -0.564283569548442
Gyc1_477 y1 0 x477 0 -0.144316333873688
Gyc1_478 y1 0 x478 0 -0.538497826265729
Gyc1_479 y1 0 x479 0 -0.093718852428342
Gyc1_480 y1 0 x480 0 0.0061847928240374
Gyc1_481 y1 0 x481 0 -0.480420484243682
Gyc1_482 y1 0 x482 0 -0.147932837565648
Gyc1_483 y1 0 x483 0 -0.555978183168216
Gyc1_484 y1 0 x484 0 1
Gyc1_485 y1 0 x485 0 -0.0162876415353556
Gyc1_486 y1 0 x486 0 0.383098873621679
Gyc1_487 y1 0 x487 0 -0.337397369338036
Gyc1_488 y1 0 x488 0 -0.730490086838918
Gyc1_489 y1 0 x489 0 -0.421920123796852
Gyc1_490 y1 0 x490 0 -0.00327605129259767
Gyc1_491 y1 0 x491 0 0.14791311656919
Gyc1_492 y1 0 x492 0 -0.110451890757927
Gyc1_493 y1 0 x493 0 -0.0232123103697893
Gyc1_494 y1 0 x494 0 -1
Gyc1_495 y1 0 x495 0 -0.109587446487652
Gyc1_496 y1 0 x496 0 0.0435371038034068
Gyc1_497 y1 0 x497 0 0.790147917097882
Gyc1_498 y1 0 x498 0 -0.104651198364276
Gyc1_499 y1 0 x499 0 -0.549792768585298
Gyc1_500 y1 0 x500 0 -0.0216563454627804
Gyc1_501 y1 0 x501 0 0.341270374022912
Gyc1_502 y1 0 x502 0 0.0271313897286925
Gyc1_503 y1 0 x503 0 0.0594998370059855
Gyc1_504 y1 0 x504 0 -0.278555738931003
Gyc1_505 y1 0 x505 0 0.10787626009938
Gyc1_506 y1 0 x506 0 0.0650629369453862
Gyc1_507 y1 0 x507 0 -0.576807908516383
Gyc1_508 y1 0 x508 0 -0.00532265685196578
Gyc1_509 y1 0 x509 0 0.883039071316271
Gyc1_510 y1 0 x510 0 -0.0676069222184878
Gyc1_511 y1 0 x511 0 -0.189899974565646
Gyc1_512 y1 0 x512 0 0.099090646023709
Gyc1_513 y1 0 x513 0 0.0185731471541693
Gyc1_514 y1 0 x514 0 0.229828443464187
Gyc1_515 y1 0 x515 0 0.0556011699261218
Gyc1_516 y1 0 x516 0 -0.0251173203640028
Gyc1_517 y1 0 x517 0 -0.0125456069625423
Gyc1_518 y1 0 x518 0 0.00493661153625739
Gyc1_519 y1 0 x519 0 0.249541279834178
Gyc1_520 y1 0 x520 0 -0.0769264144368862
Gyc1_521 y1 0 x521 0 0.0569887699804606
Gyc1_522 y1 0 x522 0 -0.0114504690420823
Gyc1_523 y1 0 x523 0 0.244416415387365
Gyc1_524 y1 0 x524 0 0.0299085037476229
Gyc1_525 y1 0 x525 0 0.0998047677141892
Gyc1_526 y1 0 x526 0 -0.159516824803057
Gyc1_527 y1 0 x527 0 0.206532616286057
Gyc1_528 y1 0 x528 0 -0.0726005638326056
Gyc1_529 y1 0 x529 0 -0.317403587052926
Gyc1_530 y1 0 x530 0 0.0424445744059234
Gyc1_531 y1 0 x531 0 -0.0675144356182053
Gyc1_532 y1 0 x532 0 -0.191128481951169
Gyc1_533 y1 0 x533 0 0.0278547358092474
Gyc1_534 y1 0 x534 0 -0.0193740620648253
Gyc1_535 y1 0 x535 0 -0.0258710537921187
Gyc1_536 y1 0 x536 0 -0.0353296791794951
Gyc1_537 y1 0 x537 0 0.0956281057305498
Gyc1_538 y1 0 x538 0 -0.0126301717570891
Gyc1_539 y1 0 x539 0 -0.00302873687695554
Gyc1_540 y1 0 x540 0 -0.195879816741542
Gyc1_541 y1 0 x541 0 0.0169759694264142
Gyc1_542 y1 0 x542 0 -0.108816569940755
Gyc1_543 y1 0 x543 0 0.0477508898502118
Gyc1_544 y1 0 x544 0 0.0281234418631045
Gyc1_545 y1 0 x545 0 0.0369393143288769
Gyc1_546 y1 0 x546 0 -0.020108859043654
Gyc1_547 y1 0 x547 0 0.0349397319160116
Gyc1_548 y1 0 x548 0 0.0461154913590748
Gyc1_549 y1 0 x549 0 -0.00826926218899498
Gyc1_550 y1 0 x550 0 -0.0938131291242225
Gyc1_551 y1 0 x551 0 -0.0249162209875939
Gyc1_552 y1 0 x552 0 -0.435020884828965
Gyc1_553 y1 0 x553 0 0.023003660850906
Gyc1_554 y1 0 x554 0 0.015031044223591
Gyc1_555 y1 0 x555 0 0.030496382371097
Gyc1_556 y1 0 x556 0 0.0813454369773643
Gyc1_557 y1 0 x557 0 0.179415221426998
Gyc1_558 y1 0 x558 0 0.278468731985576
Gyc1_559 y1 0 x559 0 0.0316428259208764
Gyc1_560 y1 0 x560 0 0.129136466637983
Gyc1_561 y1 0 x561 0 -0.00290513567462484
Gyc1_562 y1 0 x562 0 0.0600687947453261
Gyc1_563 y1 0 x563 0 0.0610491063248839
Gyc1_564 y1 0 x564 0 -0.102487564710914
Gyc1_565 y1 0 x565 0 -0.0102823281150059
Gyc1_566 y1 0 x566 0 0.0677976094660167
Gyc1_567 y1 0 x567 0 0.0416714298573413
Gyc1_568 y1 0 x568 0 0.0449444179149425
Gyc1_569 y1 0 x569 0 0.193655552182545
Gyc1_570 y1 0 x570 0 -0.0426863404856826
Gyc1_571 y1 0 x571 0 0.106819944390941
Gyc1_572 y1 0 x572 0 0.113564808586745
Gyc1_573 y1 0 x573 0 -0.0405918279497362
Gyc1_574 y1 0 x574 0 0.0194499295343392
Gyc1_575 y1 0 x575 0 0.311533254077407
Gyc1_576 y1 0 x576 0 0.0234754103004859
Gyc1_577 y1 0 x577 0 -0.107855683147564
Gyc1_578 y1 0 x578 0 0.040217067482713
Gyc1_579 y1 0 x579 0 0.127189160566792
Gyc1_580 y1 0 x580 0 0.0493923067171295
Gyc1_581 y1 0 x581 0 0.165895603379315
Gyc1_582 y1 0 x582 0 -0.0784915246184411
Gyc1_583 y1 0 x583 0 0.0683757946128622
Gyc1_584 y1 0 x584 0 -0.0267020436574554
Gyc1_585 y1 0 x585 0 0.0167278227965595
Gyc1_586 y1 0 x586 0 -0.233294463811399
Gyc1_587 y1 0 x587 0 -0.0383261195223858
Gyc1_588 y1 0 x588 0 -0.0731484154542331
Gyc1_589 y1 0 x589 0 0.0809294890041484
Gyc1_590 y1 0 x590 0 -0.104266806076306
Gyc1_591 y1 0 x591 0 -0.0801434248183695
Gyc1_592 y1 0 x592 0 0.102430407729267
Gyc1_593 y1 0 x593 0 -0.238275094483689
Gyc1_594 y1 0 x594 0 0.113836421390087
Gyc1_595 y1 0 x595 0 0.0122577237183183
Gyc1_596 y1 0 x596 0 -0.0441070356175825
Gyc1_597 y1 0 x597 0 -0.302703831563675
Gyc1_598 y1 0 x598 0 -0.293270191683904
Gyc1_599 y1 0 x599 0 -0.568630970913518
Gyc1_600 y1 0 x600 0 -0.250115389654918
Gyd1_1 y1 0 u1 0 -2.86885788860264
Gyd1_2 y1 0 u2 0 0.130304486369638
Gyd1_3 y1 0 u3 0 -0.247321117726876
Gyc2_1 y2 0 x1 0 -0.0371891324347647
Gyc2_2 y2 0 x2 0 -0.114080261585662
Gyc2_3 y2 0 x3 0 0.0287803561640079
Gyc2_4 y2 0 x4 0 -0.0683002731329166
Gyc2_5 y2 0 x5 0 -0.622992219384671
Gyc2_6 y2 0 x6 0 0.0117363267654449
Gyc2_7 y2 0 x7 0 -0.0680471314599245
Gyc2_8 y2 0 x8 0 -0.00515637070351048
Gyc2_9 y2 0 x9 0 0.0129234365584362
Gyc2_10 y2 0 x10 0 0.00337172673484183
Gyc2_11 y2 0 x11 0 0.000956354388687179
Gyc2_12 y2 0 x12 0 -0.728040813172257
Gyc2_13 y2 0 x13 0 0.192200959046323
Gyc2_14 y2 0 x14 0 -0.0948649195372484
Gyc2_15 y2 0 x15 0 -0.166389190251358
Gyc2_16 y2 0 x16 0 0.147436887365644
Gyc2_17 y2 0 x17 0 0.106071969850374
Gyc2_18 y2 0 x18 0 -0.0558078844904506
Gyc2_19 y2 0 x19 0 0.0554969400943016
Gyc2_20 y2 0 x20 0 0.0188158579646996
Gyc2_21 y2 0 x21 0 -0.0589341157210942
Gyc2_22 y2 0 x22 0 0.0388581528941402
Gyc2_23 y2 0 x23 0 0.100862103919409
Gyc2_24 y2 0 x24 0 0.00240376828754905
Gyc2_25 y2 0 x25 0 0.0299437079772337
Gyc2_26 y2 0 x26 0 -0.0599183046900402
Gyc2_27 y2 0 x27 0 -0.110926407493414
Gyc2_28 y2 0 x28 0 0.156245850534792
Gyc2_29 y2 0 x29 0 -0.0438482352730577
Gyc2_30 y2 0 x30 0 -0.532028145970712
Gyc2_31 y2 0 x31 0 0.224498150972581
Gyc2_32 y2 0 x32 0 -0.0849190086664514
Gyc2_33 y2 0 x33 0 0.0553772167122758
Gyc2_34 y2 0 x34 0 -0.16377578435658
Gyc2_35 y2 0 x35 0 0.0167668725666706
Gyc2_36 y2 0 x36 0 0.0163639926907396
Gyc2_37 y2 0 x37 0 -0.659255844359734
Gyc2_38 y2 0 x38 0 -0.00505612291134093
Gyc2_39 y2 0 x39 0 -0.598720835424949
Gyc2_40 y2 0 x40 0 -0.0859676874033454
Gyc2_41 y2 0 x41 0 -0.197035903245892
Gyc2_42 y2 0 x42 0 0.711712592414105
Gyc2_43 y2 0 x43 0 -1
Gyc2_44 y2 0 x44 0 0.148812372575533
Gyc2_45 y2 0 x45 0 0.162126187595062
Gyc2_46 y2 0 x46 0 -0.0188780348827567
Gyc2_47 y2 0 x47 0 -0.227103337470415
Gyc2_48 y2 0 x48 0 -0.0399405689837684
Gyc2_49 y2 0 x49 0 -0.0370992406252198
Gyc2_50 y2 0 x50 0 0.0266183245896723
Gyc2_51 y2 0 x51 0 -0.0363142442087672
Gyc2_52 y2 0 x52 0 0.16214711038666
Gyc2_53 y2 0 x53 0 0.0379968727238681
Gyc2_54 y2 0 x54 0 0.325873222688965
Gyc2_55 y2 0 x55 0 -0.049787338050834
Gyc2_56 y2 0 x56 0 -0.0585671183983158
Gyc2_57 y2 0 x57 0 0.901032344730759
Gyc2_58 y2 0 x58 0 0.131838391937279
Gyc2_59 y2 0 x59 0 -0.303542514400585
Gyc2_60 y2 0 x60 0 -0.201977055893624
Gyc2_61 y2 0 x61 0 -0.383626199232236
Gyc2_62 y2 0 x62 0 0.173031076865887
Gyc2_63 y2 0 x63 0 0.0613827608510841
Gyc2_64 y2 0 x64 0 -0.0100045168924542
Gyc2_65 y2 0 x65 0 -1
Gyc2_66 y2 0 x66 0 0.163168187244377
Gyc2_67 y2 0 x67 0 0.00701555486043531
Gyc2_68 y2 0 x68 0 -0.144379833870579
Gyc2_69 y2 0 x69 0 0.0162360555914929
Gyc2_70 y2 0 x70 0 -0.00101764661538083
Gyc2_71 y2 0 x71 0 -0.295742225189915
Gyc2_72 y2 0 x72 0 -1
Gyc2_73 y2 0 x73 0 -0.223035388103487
Gyc2_74 y2 0 x74 0 0.0304951536727123
Gyc2_75 y2 0 x75 0 0.200920905293714
Gyc2_76 y2 0 x76 0 -0.0863021135803506
Gyc2_77 y2 0 x77 0 -0.0630343181333981
Gyc2_78 y2 0 x78 0 -0.380815749317174
Gyc2_79 y2 0 x79 0 -0.0475931012039533
Gyc2_80 y2 0 x80 0 0.017967896641408
Gyc2_81 y2 0 x81 0 -0.992576601439924
Gyc2_82 y2 0 x82 0 -0.0546624714542453
Gyc2_83 y2 0 x83 0 -0.124803523129576
Gyc2_84 y2 0 x84 0 1
Gyc2_85 y2 0 x85 0 1
Gyc2_86 y2 0 x86 0 0.287091074553494
Gyc2_87 y2 0 x87 0 -0.291080765604271
Gyc2_88 y2 0 x88 0 -0.235407458192771
Gyc2_89 y2 0 x89 0 -0.0693859339728518
Gyc2_90 y2 0 x90 0 0.124846757103884
Gyc2_91 y2 0 x91 0 0.0203168324826294
Gyc2_92 y2 0 x92 0 -0.132607052541292
Gyc2_93 y2 0 x93 0 -0.181766768314532
Gyc2_94 y2 0 x94 0 -0.702599468773408
Gyc2_95 y2 0 x95 0 -0.450916488858369
Gyc2_96 y2 0 x96 0 0.0891759529368616
Gyc2_97 y2 0 x97 0 1
Gyc2_98 y2 0 x98 0 -0.244706789247557
Gyc2_99 y2 0 x99 0 -0.134515962882636
Gyc2_100 y2 0 x100 0 0.0509520106857484
Gyc2_101 y2 0 x101 0 0.201651516855046
Gyc2_102 y2 0 x102 0 -0.232857574646655
Gyc2_103 y2 0 x103 0 -0.167119438504001
Gyc2_104 y2 0 x104 0 -1
Gyc2_105 y2 0 x105 0 0.220474144233868
Gyc2_106 y2 0 x106 0 0.00165143340069632
Gyc2_107 y2 0 x107 0 -0.0523105328682777
Gyc2_108 y2 0 x108 0 0.659410848550316
Gyc2_109 y2 0 x109 0 0.107734789205129
Gyc2_110 y2 0 x110 0 -0.132844550919811
Gyc2_111 y2 0 x111 0 -0.152024181820267
Gyc2_112 y2 0 x112 0 0.440690936567726
Gyc2_113 y2 0 x113 0 0.0286605444200393
Gyc2_114 y2 0 x114 0 0.129935988065985
Gyc2_115 y2 0 x115 0 0.0116313215764478
Gyc2_116 y2 0 x116 0 -0.225653842514873
Gyc2_117 y2 0 x117 0 -0.0699385261613919
Gyc2_118 y2 0 x118 0 0.0156344765147724
Gyc2_119 y2 0 x119 0 0.0182774845873032
Gyc2_120 y2 0 x120 0 0.509012518469234
Gyc2_121 y2 0 x121 0 -0.0448180124980789
Gyc2_122 y2 0 x122 0 -0.0183408686490033
Gyc2_123 y2 0 x123 0 -0.00313190005702473
Gyc2_124 y2 0 x124 0 0.0210149650119193
Gyc2_125 y2 0 x125 0 -0.00877275556871401
Gyc2_126 y2 0 x126 0 0.0271872710675041
Gyc2_127 y2 0 x127 0 0.363321758466937
Gyc2_128 y2 0 x128 0 -0.315894897165232
Gyc2_129 y2 0 x129 0 -0.0294264083478889
Gyc2_130 y2 0 x130 0 -0.047671425229973
Gyc2_131 y2 0 x131 0 0.00610891958898299
Gyc2_132 y2 0 x132 0 -0.0172733912341665
Gyc2_133 y2 0 x133 0 0.0155220155355401
Gyc2_134 y2 0 x134 0 -0.0268055837203833
Gyc2_135 y2 0 x135 0 0.0141328175252574
Gyc2_136 y2 0 x136 0 -0.222080036829526
Gyc2_137 y2 0 x137 0 0.0862073459102854
Gyc2_138 y2 0 x138 0 0.0156097514301378
Gyc2_139 y2 0 x139 0 -7.91516497048087e-05
Gyc2_140 y2 0 x140 0 -0.48974737955199
Gyc2_141 y2 0 x141 0 -0.0332886412322061
Gyc2_142 y2 0 x142 0 -0.0192840448434093
Gyc2_143 y2 0 x143 0 0.0158116071705226
Gyc2_144 y2 0 x144 0 -0.0500525380101617
Gyc2_145 y2 0 x145 0 0.0744541182694807
Gyc2_146 y2 0 x146 0 -0.081872709901986
Gyc2_147 y2 0 x147 0 0.0559145964004257
Gyc2_148 y2 0 x148 0 0.216169900395539
Gyc2_149 y2 0 x149 0 0.0503313314505329
Gyc2_150 y2 0 x150 0 -0.471665242994545
Gyc2_151 y2 0 x151 0 -0.0135546335521752
Gyc2_152 y2 0 x152 0 -0.179164773693493
Gyc2_153 y2 0 x153 0 0.0226716639776931
Gyc2_154 y2 0 x154 0 -0.0498240931526031
Gyc2_155 y2 0 x155 0 -0.216715886007105
Gyc2_156 y2 0 x156 0 0.0471020151363368
Gyc2_157 y2 0 x157 0 0.657645233699375
Gyc2_158 y2 0 x158 0 -0.00944889900210701
Gyc2_159 y2 0 x159 0 0.0842139836958434
Gyc2_160 y2 0 x160 0 -0.00641185846363823
Gyc2_161 y2 0 x161 0 0.0314280813113574
Gyc2_162 y2 0 x162 0 -0.00103829520768918
Gyc2_163 y2 0 x163 0 0.0629664125415677
Gyc2_164 y2 0 x164 0 -0.0541813584932864
Gyc2_165 y2 0 x165 0 -0.147555732874196
Gyc2_166 y2 0 x166 0 -0.031166699772268
Gyc2_167 y2 0 x167 0 -0.0525605977459975
Gyc2_168 y2 0 x168 0 -0.0404350757843722
Gyc2_169 y2 0 x169 0 0.235855610038194
Gyc2_170 y2 0 x170 0 0.0505976287742434
Gyc2_171 y2 0 x171 0 0.226532052738668
Gyc2_172 y2 0 x172 0 0.0343917681043389
Gyc2_173 y2 0 x173 0 0.00314312200304228
Gyc2_174 y2 0 x174 0 -0.0504429614901966
Gyc2_175 y2 0 x175 0 0.251345940825075
Gyc2_176 y2 0 x176 0 0.110575960752996
Gyc2_177 y2 0 x177 0 0.0506999281059677
Gyc2_178 y2 0 x178 0 -0.0205327874080288
Gyc2_179 y2 0 x179 0 0.403378858787944
Gyc2_180 y2 0 x180 0 0.00318955915445481
Gyc2_181 y2 0 x181 0 0.0586161503544318
Gyc2_182 y2 0 x182 0 0.00363290785913551
Gyc2_183 y2 0 x183 0 0.0299566308625526
Gyc2_184 y2 0 x184 0 0.0645803993200554
Gyc2_185 y2 0 x185 0 0.103206162941227
Gyc2_186 y2 0 x186 0 -0.12420212985942
Gyc2_187 y2 0 x187 0 0.0950898740541416
Gyc2_188 y2 0 x188 0 0.0264537056548608
Gyc2_189 y2 0 x189 0 0.00447458434062156
Gyc2_190 y2 0 x190 0 0.155565444931455
Gyc2_191 y2 0 x191 0 -0.00802339655771713
Gyc2_192 y2 0 x192 0 -0.124803639269588
Gyc2_193 y2 0 x193 0 0.0604855306276694
Gyc2_194 y2 0 x194 0 0.0212513552238404
Gyc2_195 y2 0 x195 0 -0.012332773970685
Gyc2_196 y2 0 x196 0 -0.00464257797444241
Gyc2_197 y2 0 x197 0 0.0814563901227946
Gyc2_198 y2 0 x198 0 0.1641113314055
Gyc2_199 y2 0 x199 0 0.526805297481526
Gyc2_200 y2 0 x200 0 0.453625944739642
Gyc2_201 y2 0 x201 0 -0.803233144346733
Gyc2_202 y2 0 x202 0 1
Gyc2_203 y2 0 x203 0 1
Gyc2_204 y2 0 x204 0 1
Gyc2_205 y2 0 x205 0 1
Gyc2_206 y2 0 x206 0 1
Gyc2_207 y2 0 x207 0 -1
Gyc2_208 y2 0 x208 0 1
Gyc2_209 y2 0 x209 0 -1
Gyc2_210 y2 0 x210 0 0.777627609927711
Gyc2_211 y2 0 x211 0 -1
Gyc2_212 y2 0 x212 0 1
Gyc2_213 y2 0 x213 0 -1
Gyc2_214 y2 0 x214 0 -0.677562657192568
Gyc2_215 y2 0 x215 0 -0.797627563539484
Gyc2_216 y2 0 x216 0 -1
Gyc2_217 y2 0 x217 0 0.153219098653993
Gyc2_218 y2 0 x218 0 -1
Gyc2_219 y2 0 x219 0 1
Gyc2_220 y2 0 x220 0 -1
Gyc2_221 y2 0 x221 0 1
Gyc2_222 y2 0 x222 0 -0.604026814992313
Gyc2_223 y2 0 x223 0 1
Gyc2_224 y2 0 x224 0 1
Gyc2_225 y2 0 x225 0 1
Gyc2_226 y2 0 x226 0 0.67842422423842
Gyc2_227 y2 0 x227 0 -0.792189900132051
Gyc2_228 y2 0 x228 0 -1
Gyc2_229 y2 0 x229 0 -0.714933207338573
Gyc2_230 y2 0 x230 0 0.258569941638594
Gyc2_231 y2 0 x231 0 -1
Gyc2_232 y2 0 x232 0 -0.721381767151298
Gyc2_233 y2 0 x233 0 1
Gyc2_234 y2 0 x234 0 -1
Gyc2_235 y2 0 x235 0 -1
Gyc2_236 y2 0 x236 0 -1
Gyc2_237 y2 0 x237 0 0.58735431462316
Gyc2_238 y2 0 x238 0 0.75658664075099
Gyc2_239 y2 0 x239 0 -1
Gyc2_240 y2 0 x240 0 -1
Gyc2_241 y2 0 x241 0 -0.242001856122801
Gyc2_242 y2 0 x242 0 -0.669092101300215
Gyc2_243 y2 0 x243 0 0.407574934840992
Gyc2_244 y2 0 x244 0 0.723467281381648
Gyc2_245 y2 0 x245 0 1
Gyc2_246 y2 0 x246 0 0.371190369182656
Gyc2_247 y2 0 x247 0 0.0959868103305968
Gyc2_248 y2 0 x248 0 -0.867086896969184
Gyc2_249 y2 0 x249 0 0.990948367980017
Gyc2_250 y2 0 x250 0 0.534277095744391
Gyc2_251 y2 0 x251 0 1
Gyc2_252 y2 0 x252 0 1
Gyc2_253 y2 0 x253 0 -0.65091786341863
Gyc2_254 y2 0 x254 0 0.774036834553658
Gyc2_255 y2 0 x255 0 0.249512536912514
Gyc2_256 y2 0 x256 0 0.601357085438662
Gyc2_257 y2 0 x257 0 -0.342342792569971
Gyc2_258 y2 0 x258 0 -0.0352737796230673
Gyc2_259 y2 0 x259 0 -0.481455921124742
Gyc2_260 y2 0 x260 0 1
Gyc2_261 y2 0 x261 0 -0.526597304192434
Gyc2_262 y2 0 x262 0 1
Gyc2_263 y2 0 x263 0 -0.440326331023922
Gyc2_264 y2 0 x264 0 0.55287027105284
Gyc2_265 y2 0 x265 0 0.091624867623034
Gyc2_266 y2 0 x266 0 1
Gyc2_267 y2 0 x267 0 1
Gyc2_268 y2 0 x268 0 0.189857764158707
Gyc2_269 y2 0 x269 0 -0.0753048684927983
Gyc2_270 y2 0 x270 0 1
Gyc2_271 y2 0 x271 0 -1
Gyc2_272 y2 0 x272 0 1
Gyc2_273 y2 0 x273 0 -1
Gyc2_274 y2 0 x274 0 1
Gyc2_275 y2 0 x275 0 -0.00254334952451899
Gyc2_276 y2 0 x276 0 -0.664595686095802
Gyc2_277 y2 0 x277 0 -1
Gyc2_278 y2 0 x278 0 -1
Gyc2_279 y2 0 x279 0 -0.500316922643513
Gyc2_280 y2 0 x280 0 0.391175426088777
Gyc2_281 y2 0 x281 0 -0.555456840656911
Gyc2_282 y2 0 x282 0 0.411477202961145
Gyc2_283 y2 0 x283 0 0.0859786047458894
Gyc2_284 y2 0 x284 0 1
Gyc2_285 y2 0 x285 0 1
Gyc2_286 y2 0 x286 0 -0.0532428375173779
Gyc2_287 y2 0 x287 0 -0.847545098863666
Gyc2_288 y2 0 x288 0 -0.0584214487884198
Gyc2_289 y2 0 x289 0 0.492517118407421
Gyc2_290 y2 0 x290 0 0.296094510132405
Gyc2_291 y2 0 x291 0 1
Gyc2_292 y2 0 x292 0 -1
Gyc2_293 y2 0 x293 0 -0.877625588509596
Gyc2_294 y2 0 x294 0 -0.29135303947786
Gyc2_295 y2 0 x295 0 1
Gyc2_296 y2 0 x296 0 1
Gyc2_297 y2 0 x297 0 0.492936981118714
Gyc2_298 y2 0 x298 0 -0.226435032921762
Gyc2_299 y2 0 x299 0 0.9203263579263
Gyc2_300 y2 0 x300 0 1
Gyc2_301 y2 0 x301 0 0.535059245367985
Gyc2_302 y2 0 x302 0 0.346602482258871
Gyc2_303 y2 0 x303 0 0.0988574505282798
Gyc2_304 y2 0 x304 0 0.458822096955636
Gyc2_305 y2 0 x305 0 1
Gyc2_306 y2 0 x306 0 -1
Gyc2_307 y2 0 x307 0 0.64235776015513
Gyc2_308 y2 0 x308 0 1
Gyc2_309 y2 0 x309 0 -0.510678156718128
Gyc2_310 y2 0 x310 0 -1
Gyc2_311 y2 0 x311 0 0.12267126182343
Gyc2_312 y2 0 x312 0 -0.582887997475626
Gyc2_313 y2 0 x313 0 0.436879896588105
Gyc2_314 y2 0 x314 0 0.231994225678199
Gyc2_315 y2 0 x315 0 -1
Gyc2_316 y2 0 x316 0 1
Gyc2_317 y2 0 x317 0 1
Gyc2_318 y2 0 x318 0 1
Gyc2_319 y2 0 x319 0 -1
Gyc2_320 y2 0 x320 0 0.727337207741572
Gyc2_321 y2 0 x321 0 0.173274608864607
Gyc2_322 y2 0 x322 0 1
Gyc2_323 y2 0 x323 0 -0.593346099789435
Gyc2_324 y2 0 x324 0 0.841855168521206
Gyc2_325 y2 0 x325 0 -0.248566446912124
Gyc2_326 y2 0 x326 0 0.608659822811247
Gyc2_327 y2 0 x327 0 0.562005317659806
Gyc2_328 y2 0 x328 0 -1
Gyc2_329 y2 0 x329 0 0.69156653309448
Gyc2_330 y2 0 x330 0 -1
Gyc2_331 y2 0 x331 0 -0.152662660926124
Gyc2_332 y2 0 x332 0 0.197533036240107
Gyc2_333 y2 0 x333 0 1
Gyc2_334 y2 0 x334 0 -0.084792140056974
Gyc2_335 y2 0 x335 0 -1
Gyc2_336 y2 0 x336 0 1
Gyc2_337 y2 0 x337 0 0.0755181555373763
Gyc2_338 y2 0 x338 0 0.316505534885078
Gyc2_339 y2 0 x339 0 1
Gyc2_340 y2 0 x340 0 0.701477974412731
Gyc2_341 y2 0 x341 0 0.38237115372477
Gyc2_342 y2 0 x342 0 0.396091735791118
Gyc2_343 y2 0 x343 0 1
Gyc2_344 y2 0 x344 0 0.0360034169160282
Gyc2_345 y2 0 x345 0 -0.707140145872763
Gyc2_346 y2 0 x346 0 0.317392657179271
Gyc2_347 y2 0 x347 0 1
Gyc2_348 y2 0 x348 0 -1
Gyc2_349 y2 0 x349 0 -0.0458413786076003
Gyc2_350 y2 0 x350 0 -0.660625760020697
Gyc2_351 y2 0 x351 0 0.885582006852881
Gyc2_352 y2 0 x352 0 1
Gyc2_353 y2 0 x353 0 0.019476720922911
Gyc2_354 y2 0 x354 0 -1
Gyc2_355 y2 0 x355 0 -1
Gyc2_356 y2 0 x356 0 -0.517490772977341
Gyc2_357 y2 0 x357 0 -1
Gyc2_358 y2 0 x358 0 0.341629509752524
Gyc2_359 y2 0 x359 0 -0.588621162932042
Gyc2_360 y2 0 x360 0 -0.238154181724531
Gyc2_361 y2 0 x361 0 -0.304127485833164
Gyc2_362 y2 0 x362 0 0.143795817003785
Gyc2_363 y2 0 x363 0 -0.499719455970658
Gyc2_364 y2 0 x364 0 -0.327421908217518
Gyc2_365 y2 0 x365 0 0.731973147909612
Gyc2_366 y2 0 x366 0 0.18570179310699
Gyc2_367 y2 0 x367 0 1
Gyc2_368 y2 0 x368 0 0.0973044652266858
Gyc2_369 y2 0 x369 0 -0.869877668218608
Gyc2_370 y2 0 x370 0 -0.344083107602237
Gyc2_371 y2 0 x371 0 1
Gyc2_372 y2 0 x372 0 -0.0803431441801868
Gyc2_373 y2 0 x373 0 0.101726603519895
Gyc2_374 y2 0 x374 0 0.489383352848709
Gyc2_375 y2 0 x375 0 -0.252297116556349
Gyc2_376 y2 0 x376 0 -0.372279231494473
Gyc2_377 y2 0 x377 0 -0.145966367315274
Gyc2_378 y2 0 x378 0 0.134013531230076
Gyc2_379 y2 0 x379 0 0.535639697370792
Gyc2_380 y2 0 x380 0 -0.0283214529117885
Gyc2_381 y2 0 x381 0 -0.247999373315412
Gyc2_382 y2 0 x382 0 0.138240068625109
Gyc2_383 y2 0 x383 0 -0.358093642362964
Gyc2_384 y2 0 x384 0 -0.748013795144143
Gyc2_385 y2 0 x385 0 -0.564980233876798
Gyc2_386 y2 0 x386 0 0.329390531184792
Gyc2_387 y2 0 x387 0 -1
Gyc2_388 y2 0 x388 0 0.0626354860565176
Gyc2_389 y2 0 x389 0 -0.194660997542055
Gyc2_390 y2 0 x390 0 -0.989472856908032
Gyc2_391 y2 0 x391 0 0.214778887582962
Gyc2_392 y2 0 x392 0 0.949028886364576
Gyc2_393 y2 0 x393 0 0.620819593270959
Gyc2_394 y2 0 x394 0 0.11331490790109
Gyc2_395 y2 0 x395 0 1
Gyc2_396 y2 0 x396 0 0.164596270044907
Gyc2_397 y2 0 x397 0 -0.116626608228226
Gyc2_398 y2 0 x398 0 -0.31201949889461
Gyc2_399 y2 0 x399 0 1
Gyc2_400 y2 0 x400 0 1
Gyc2_401 y2 0 x401 0 -0.263361890084449
Gyc2_402 y2 0 x402 0 0.112675097135364
Gyc2_403 y2 0 x403 0 -0.111444153468536
Gyc2_404 y2 0 x404 0 0.166674152599354
Gyc2_405 y2 0 x405 0 -0.0764388623517309
Gyc2_406 y2 0 x406 0 0.203077100422084
Gyc2_407 y2 0 x407 0 -1
Gyc2_408 y2 0 x408 0 0.0105356855784979
Gyc2_409 y2 0 x409 0 -0.0692134292660573
Gyc2_410 y2 0 x410 0 -0.277401442283861
Gyc2_411 y2 0 x411 0 -0.266275420390129
Gyc2_412 y2 0 x412 0 -0.0562110704089811
Gyc2_413 y2 0 x413 0 -0.075326925255027
Gyc2_414 y2 0 x414 0 -0.823870063468276
Gyc2_415 y2 0 x415 0 0.364233716570468
Gyc2_416 y2 0 x416 0 0.0468534581865577
Gyc2_417 y2 0 x417 0 0.925079096635363
Gyc2_418 y2 0 x418 0 -0.206113765068829
Gyc2_419 y2 0 x419 0 0.272973799162744
Gyc2_420 y2 0 x420 0 0.00540488712128529
Gyc2_421 y2 0 x421 0 0.0377440241483645
Gyc2_422 y2 0 x422 0 0.707082713524124
Gyc2_423 y2 0 x423 0 0.0123374065574441
Gyc2_424 y2 0 x424 0 0.246105023948673
Gyc2_425 y2 0 x425 0 -0.0367259473544177
Gyc2_426 y2 0 x426 0 0.215731651076886
Gyc2_427 y2 0 x427 0 0.353293689614233
Gyc2_428 y2 0 x428 0 -0.0510295473167127
Gyc2_429 y2 0 x429 0 -0.848295313626674
Gyc2_430 y2 0 x430 0 -0.0257044134134758
Gyc2_431 y2 0 x431 0 0.000249124997141201
Gyc2_432 y2 0 x432 0 -0.58122218443774
Gyc2_433 y2 0 x433 0 0.316222326697894
Gyc2_434 y2 0 x434 0 0.112366827736396
Gyc2_435 y2 0 x435 0 0.326644428660088
Gyc2_436 y2 0 x436 0 -0.203794852045612
Gyc2_437 y2 0 x437 0 -0.0604267125440127
Gyc2_438 y2 0 x438 0 0.345278471456607
Gyc2_439 y2 0 x439 0 0.197448338899691
Gyc2_440 y2 0 x440 0 -0.274123659487098
Gyc2_441 y2 0 x441 0 0.571363167485269
Gyc2_442 y2 0 x442 0 -0.0136545660839444
Gyc2_443 y2 0 x443 0 0.0674403816614329
Gyc2_444 y2 0 x444 0 0.79280504197231
Gyc2_445 y2 0 x445 0 -0.00281170592960444
Gyc2_446 y2 0 x446 0 0.362826591330452
Gyc2_447 y2 0 x447 0 0.178728224456101
Gyc2_448 y2 0 x448 0 0.3019806611082
Gyc2_449 y2 0 x449 0 0.167863357964165
Gyc2_450 y2 0 x450 0 0.265655517721297
Gyc2_451 y2 0 x451 0 -0.629709885423552
Gyc2_452 y2 0 x452 0 0.249284216532051
Gyc2_453 y2 0 x453 0 -0.121393515702085
Gyc2_454 y2 0 x454 0 -0.658143221119908
Gyc2_455 y2 0 x455 0 -1
Gyc2_456 y2 0 x456 0 0.26007626259545
Gyc2_457 y2 0 x457 0 0.0340958859123738
Gyc2_458 y2 0 x458 0 -0.456912475841783
Gyc2_459 y2 0 x459 0 -0.592475477081293
Gyc2_460 y2 0 x460 0 -1
Gyc2_461 y2 0 x461 0 0.229549968045526
Gyc2_462 y2 0 x462 0 0.0597053918282838
Gyc2_463 y2 0 x463 0 -0.271316705984181
Gyc2_464 y2 0 x464 0 -1
Gyc2_465 y2 0 x465 0 0.0395407501399135
Gyc2_466 y2 0 x466 0 0.976861740317166
Gyc2_467 y2 0 x467 0 0.145709651952634
Gyc2_468 y2 0 x468 0 0.251241519862794
Gyc2_469 y2 0 x469 0 -0.517159653579119
Gyc2_470 y2 0 x470 0 0.151318619713597
Gyc2_471 y2 0 x471 0 -0.55865644597908
Gyc2_472 y2 0 x472 0 0.173212361206896
Gyc2_473 y2 0 x473 0 -0.400493940324973
Gyc2_474 y2 0 x474 0 0.0081824773258027
Gyc2_475 y2 0 x475 0 -0.225585306981522
Gyc2_476 y2 0 x476 0 -0.469107185167129
Gyc2_477 y2 0 x477 0 0.180478670924855
Gyc2_478 y2 0 x478 0 -0.411224887636784
Gyc2_479 y2 0 x479 0 -0.35471160647739
Gyc2_480 y2 0 x480 0 -0.361860050026254
Gyc2_481 y2 0 x481 0 -0.0164493085011205
Gyc2_482 y2 0 x482 0 0.555576389589427
Gyc2_483 y2 0 x483 0 -0.466248812027914
Gyc2_484 y2 0 x484 0 0.79662793565649
Gyc2_485 y2 0 x485 0 -0.0140781912597531
Gyc2_486 y2 0 x486 0 -0.280028550092735
Gyc2_487 y2 0 x487 0 0.259477334309415
Gyc2_488 y2 0 x488 0 -0.535964524191361
Gyc2_489 y2 0 x489 0 0.504996921492952
Gyc2_490 y2 0 x490 0 -0.418458553874203
Gyc2_491 y2 0 x491 0 0.0219492515831927
Gyc2_492 y2 0 x492 0 -0.121026551549825
Gyc2_493 y2 0 x493 0 0.33770406314864
Gyc2_494 y2 0 x494 0 0.299464813435762
Gyc2_495 y2 0 x495 0 0.076536438279926
Gyc2_496 y2 0 x496 0 0.0138177980892159
Gyc2_497 y2 0 x497 0 -0.538590560786593
Gyc2_498 y2 0 x498 0 0.271845155151757
Gyc2_499 y2 0 x499 0 -0.628821989053806
Gyc2_500 y2 0 x500 0 0.0675506580987192
Gyc2_501 y2 0 x501 0 -1
Gyc2_502 y2 0 x502 0 0.157444651303333
Gyc2_503 y2 0 x503 0 -1
Gyc2_504 y2 0 x504 0 0.345257709777796
Gyc2_505 y2 0 x505 0 -0.15137654159944
Gyc2_506 y2 0 x506 0 -0.0736594209352693
Gyc2_507 y2 0 x507 0 -0.854809877172298
Gyc2_508 y2 0 x508 0 -0.202107189327131
Gyc2_509 y2 0 x509 0 1
Gyc2_510 y2 0 x510 0 -0.21928622225821
Gyc2_511 y2 0 x511 0 0.92176680517617
Gyc2_512 y2 0 x512 0 -0.080426535657883
Gyc2_513 y2 0 x513 0 0.337535712197284
Gyc2_514 y2 0 x514 0 0.448678514261286
Gyc2_515 y2 0 x515 0 -0.218396941275825
Gyc2_516 y2 0 x516 0 -0.0983736140143899
Gyc2_517 y2 0 x517 0 0.139243626644858
Gyc2_518 y2 0 x518 0 0.182841887099068
Gyc2_519 y2 0 x519 0 0.844283298858767
Gyc2_520 y2 0 x520 0 -0.711461631346841
Gyc2_521 y2 0 x521 0 0.227358209694649
Gyc2_522 y2 0 x522 0 0.174483985306248
Gyc2_523 y2 0 x523 0 1
Gyc2_524 y2 0 x524 0 0.201410532530655
Gyc2_525 y2 0 x525 0 0.626814704525707
Gyc2_526 y2 0 x526 0 -0.341619598520681
Gyc2_527 y2 0 x527 0 -0.0482535465553953
Gyc2_528 y2 0 x528 0 -0.192090025994798
Gyc2_529 y2 0 x529 0 -0.715417612300148
Gyc2_530 y2 0 x530 0 0.22205046318741
Gyc2_531 y2 0 x531 0 -0.383870170785407
Gyc2_532 y2 0 x532 0 -0.654042978388811
Gyc2_533 y2 0 x533 0 0.192386611699068
Gyc2_534 y2 0 x534 0 0.632851365348486
Gyc2_535 y2 0 x535 0 -0.00253643158339097
Gyc2_536 y2 0 x536 0 0.161397461229024
Gyc2_537 y2 0 x537 0 0.773249274625264
Gyc2_538 y2 0 x538 0 -0.746789169733163
Gyc2_539 y2 0 x539 0 0.114210758148228
Gyc2_540 y2 0 x540 0 -1
Gyc2_541 y2 0 x541 0 0.43150122492105
Gyc2_542 y2 0 x542 0 -0.84043578513836
Gyc2_543 y2 0 x543 0 0.216508635627813
Gyc2_544 y2 0 x544 0 0.939976010156425
Gyc2_545 y2 0 x545 0 -0.0627833436160021
Gyc2_546 y2 0 x546 0 -0.423185696567333
Gyc2_547 y2 0 x547 0 0.0987006468181164
Gyc2_548 y2 0 x548 0 0.137757917571267
Gyc2_549 y2 0 x549 0 -0.568576542602185
Gyc2_550 y2 0 x550 0 -0.187854527478776
Gyc2_551 y2 0 x551 0 -0.62898521113685
Gyc2_552 y2 0 x552 0 0.325416364704548
Gyc2_553 y2 0 x553 0 -0.357752519116938
Gyc2_554 y2 0 x554 0 0.0368990081816535
Gyc2_555 y2 0 x555 0 0.282725960200733
Gyc2_556 y2 0 x556 0 -0.233361493651029
Gyc2_557 y2 0 x557 0 -0.134971480803137
Gyc2_558 y2 0 x558 0 1
Gyc2_559 y2 0 x559 0 -0.342106410377639
Gyc2_560 y2 0 x560 0 1
Gyc2_561 y2 0 x561 0 -0.362423983568056
Gyc2_562 y2 0 x562 0 -0.720702356471066
Gyc2_563 y2 0 x563 0 0.44014957465333
Gyc2_564 y2 0 x564 0 -0.300803003835702
Gyc2_565 y2 0 x565 0 0.373833575715367
Gyc2_566 y2 0 x566 0 0.785583475596483
Gyc2_567 y2 0 x567 0 0.114935521697703
Gyc2_568 y2 0 x568 0 0.496250876264352
Gyc2_569 y2 0 x569 0 -0.0329083831332733
Gyc2_570 y2 0 x570 0 -0.453012096093596
Gyc2_571 y2 0 x571 0 0.0191188254057853
Gyc2_572 y2 0 x572 0 0.383485950048002
Gyc2_573 y2 0 x573 0 -0.670210540978736
Gyc2_574 y2 0 x574 0 0.293789750213956
Gyc2_575 y2 0 x575 0 0.858233337203627
Gyc2_576 y2 0 x576 0 -0.432039527819047
Gyc2_577 y2 0 x577 0 -0.27014532476152
Gyc2_578 y2 0 x578 0 -0.845239118631657
Gyc2_579 y2 0 x579 0 -0.161660922013791
Gyc2_580 y2 0 x580 0 0.373892562110196
Gyc2_581 y2 0 x581 0 0.270273286131605
Gyc2_582 y2 0 x582 0 0.541567902063428
Gyc2_583 y2 0 x583 0 0.920788779224483
Gyc2_584 y2 0 x584 0 -0.250115499486963
Gyc2_585 y2 0 x585 0 -0.392317392867026
Gyc2_586 y2 0 x586 0 -1
Gyc2_587 y2 0 x587 0 -0.0850295551748504
Gyc2_588 y2 0 x588 0 -0.609313059930721
Gyc2_589 y2 0 x589 0 0.576503359442024
Gyc2_590 y2 0 x590 0 -0.100770433020964
Gyc2_591 y2 0 x591 0 -0.608049203767101
Gyc2_592 y2 0 x592 0 0.140594539069772
Gyc2_593 y2 0 x593 0 -0.0515343191902169
Gyc2_594 y2 0 x594 0 -0.870242063993855
Gyc2_595 y2 0 x595 0 0.000244103044858497
Gyc2_596 y2 0 x596 0 0.547232217958848
Gyc2_597 y2 0 x597 0 1
Gyc2_598 y2 0 x598 0 -0.0635127041644143
Gyc2_599 y2 0 x599 0 0.568702805712523
Gyc2_600 y2 0 x600 0 0.654925090898198
Gyd2_1 y2 0 u1 0 0.149504352457505
Gyd2_2 y2 0 u2 0 -0.698387151400012
Gyd2_3 y2 0 u3 0 -0.57409102200985
Gyc3_1 y3 0 x1 0 -0.0785307083649798
Gyc3_2 y3 0 x2 0 0.139948102451112
Gyc3_3 y3 0 x3 0 -0.0349172053252227
Gyc3_4 y3 0 x4 0 0.136011132754329
Gyc3_5 y3 0 x5 0 -1
Gyc3_6 y3 0 x6 0 0.0444581217956148
Gyc3_7 y3 0 x7 0 -0.103833078879605
Gyc3_8 y3 0 x8 0 -0.151613006278156
Gyc3_9 y3 0 x9 0 0.0523600504299353
Gyc3_10 y3 0 x10 0 -0.0266562519822826
Gyc3_11 y3 0 x11 0 0.00873569050662523
Gyc3_12 y3 0 x12 0 -1
Gyc3_13 y3 0 x13 0 0.20768840866953
Gyc3_14 y3 0 x14 0 -0.123587518254425
Gyc3_15 y3 0 x15 0 0.491920700624988
Gyc3_16 y3 0 x16 0 -0.289464889059234
Gyc3_17 y3 0 x17 0 0.115820594331572
Gyc3_18 y3 0 x18 0 -0.0941936378942689
Gyc3_19 y3 0 x19 0 0.10356477252676
Gyc3_20 y3 0 x20 0 -0.016220663293856
Gyc3_21 y3 0 x21 0 -0.0022859281609752
Gyc3_22 y3 0 x22 0 0.00028505488989017
Gyc3_23 y3 0 x23 0 0.0723208508450425
Gyc3_24 y3 0 x24 0 0.0808940937099314
Gyc3_25 y3 0 x25 0 0.120963801162125
Gyc3_26 y3 0 x26 0 0.0587282946996534
Gyc3_27 y3 0 x27 0 0.021696846840797
Gyc3_28 y3 0 x28 0 -0.48088899439698
Gyc3_29 y3 0 x29 0 0.0470493228551235
Gyc3_30 y3 0 x30 0 0.11522009237002
Gyc3_31 y3 0 x31 0 0.0347361462663412
Gyc3_32 y3 0 x32 0 0.0551485288840684
Gyc3_33 y3 0 x33 0 0.00974650937509858
Gyc3_34 y3 0 x34 0 0.335889787985689
Gyc3_35 y3 0 x35 0 0.0499821832760007
Gyc3_36 y3 0 x36 0 -0.0290224667267065
Gyc3_37 y3 0 x37 0 0.224743771077058
Gyc3_38 y3 0 x38 0 0.0100307090499894
Gyc3_39 y3 0 x39 0 0.449793605760982
Gyc3_40 y3 0 x40 0 0.00966030895011428
Gyc3_41 y3 0 x41 0 0.135327057226581
Gyc3_42 y3 0 x42 0 0.1870719222405
Gyc3_43 y3 0 x43 0 0.563752562605943
Gyc3_44 y3 0 x44 0 0.0559213823800359
Gyc3_45 y3 0 x45 0 -0.407604890700199
Gyc3_46 y3 0 x46 0 0.0221822972415603
Gyc3_47 y3 0 x47 0 0.0760750132541192
Gyc3_48 y3 0 x48 0 0.28740630144434
Gyc3_49 y3 0 x49 0 0.0792172658511202
Gyc3_50 y3 0 x50 0 0.0164542568597409
Gyc3_51 y3 0 x51 0 0.12978321227907
Gyc3_52 y3 0 x52 0 0.0140172857156851
Gyc3_53 y3 0 x53 0 0.208517420768072
Gyc3_54 y3 0 x54 0 -0.129983458218631
Gyc3_55 y3 0 x55 0 -0.118010000696166
Gyc3_56 y3 0 x56 0 0.055657815765028
Gyc3_57 y3 0 x57 0 0.445589948303962
Gyc3_58 y3 0 x58 0 -0.0923942991546822
Gyc3_59 y3 0 x59 0 -0.592578743580528
Gyc3_60 y3 0 x60 0 0.0296518617569195
Gyc3_61 y3 0 x61 0 0.00690283550279565
Gyc3_62 y3 0 x62 0 1
Gyc3_63 y3 0 x63 0 -0.0756540781344204
Gyc3_64 y3 0 x64 0 -0.0399901289883987
Gyc3_65 y3 0 x65 0 -0.077365666297357
Gyc3_66 y3 0 x66 0 0.26205860685565
Gyc3_67 y3 0 x67 0 -0.0327722819016367
Gyc3_68 y3 0 x68 0 -0.0580676428914178
Gyc3_69 y3 0 x69 0 -0.0609063583914299
Gyc3_70 y3 0 x70 0 0.0394632956316072
Gyc3_71 y3 0 x71 0 -0.373590578434293
Gyc3_72 y3 0 x72 0 0.149994544525834
Gyc3_73 y3 0 x73 0 -0.240508099142688
Gyc3_74 y3 0 x74 0 0.109940953114868
Gyc3_75 y3 0 x75 0 0.128908342720262
Gyc3_76 y3 0 x76 0 -0.259618973150898
Gyc3_77 y3 0 x77 0 -0.0566886575014503
Gyc3_78 y3 0 x78 0 -0.399290841534777
Gyc3_79 y3 0 x79 0 -0.0889138680823083
Gyc3_80 y3 0 x80 0 -0.0183256193422629
Gyc3_81 y3 0 x81 0 -0.999837322514809
Gyc3_82 y3 0 x82 0 -0.0326795461527143
Gyc3_83 y3 0 x83 0 -0.200055356886704
Gyc3_84 y3 0 x84 0 0.988066549148632
Gyc3_85 y3 0 x85 0 0.143409088824313
Gyc3_86 y3 0 x86 0 0.260723050224032
Gyc3_87 y3 0 x87 0 -0.110964770531271
Gyc3_88 y3 0 x88 0 -0.314018722256854
Gyc3_89 y3 0 x89 0 -0.0987665475582068
Gyc3_90 y3 0 x90 0 -0.0266238008696404
Gyc3_91 y3 0 x91 0 0.108451758425899
Gyc3_92 y3 0 x92 0 -0.134198612888958
Gyc3_93 y3 0 x93 0 -0.011602156434307
Gyc3_94 y3 0 x94 0 -0.989422669078672
Gyc3_95 y3 0 x95 0 -0.642660498706747
Gyc3_96 y3 0 x96 0 0.0612269087325707
Gyc3_97 y3 0 x97 0 0.930265453061326
Gyc3_98 y3 0 x98 0 -0.0551486476180178
Gyc3_99 y3 0 x99 0 -0.111193289560727
Gyc3_100 y3 0 x100 0 -0.0302540335681772
Gyc3_101 y3 0 x101 0 0.101210075498737
Gyc3_102 y3 0 x102 0 0.0495503330617825
Gyc3_103 y3 0 x103 0 -0.0153912230036658
Gyc3_104 y3 0 x104 0 -0.690362411273512
Gyc3_105 y3 0 x105 0 0.0573962985035918
Gyc3_106 y3 0 x106 0 0.0500643964305141
Gyc3_107 y3 0 x107 0 -0.141874199691791
Gyc3_108 y3 0 x108 0 -0.00702207402806318
Gyc3_109 y3 0 x109 0 0.138928292565853
Gyc3_110 y3 0 x110 0 -0.0691349453968725
Gyc3_111 y3 0 x111 0 -0.0634930889876599
Gyc3_112 y3 0 x112 0 0.174243235809054
Gyc3_113 y3 0 x113 0 0.0265816767794885
Gyc3_114 y3 0 x114 0 0.0992858261149914
Gyc3_115 y3 0 x115 0 0.0995900770699359
Gyc3_116 y3 0 x116 0 -0.118126217697256
Gyc3_117 y3 0 x117 0 -0.0435948552997385
Gyc3_118 y3 0 x118 0 0.0262216304704326
Gyc3_119 y3 0 x119 0 0.0910765029521808
Gyc3_120 y3 0 x120 0 -0.0572531390774679
Gyc3_121 y3 0 x121 0 0.0342789732181171
Gyc3_122 y3 0 x122 0 0.00109630543560913
Gyc3_123 y3 0 x123 0 0.0700171091146031
Gyc3_124 y3 0 x124 0 0.0499510116444817
Gyc3_125 y3 0 x125 0 0.0439052548111515
Gyc3_126 y3 0 x126 0 -0.0502575459488559
Gyc3_127 y3 0 x127 0 0.265698676020588
Gyc3_128 y3 0 x128 0 -0.426460977644938
Gyc3_129 y3 0 x129 0 -0.0763876737814673
Gyc3_130 y3 0 x130 0 0.0620770547460875
Gyc3_131 y3 0 x131 0 -0.0552416468099251
Gyc3_132 y3 0 x132 0 -0.0922157523799206
Gyc3_133 y3 0 x133 0 0.0882779894227478
Gyc3_134 y3 0 x134 0 0.00366771696326921
Gyc3_135 y3 0 x135 0 -0.0509891841841607
Gyc3_136 y3 0 x136 0 -0.147873446971334
Gyc3_137 y3 0 x137 0 0.114930945187978
Gyc3_138 y3 0 x138 0 -0.0277795315561264
Gyc3_139 y3 0 x139 0 0.0228364303537858
Gyc3_140 y3 0 x140 0 -0.325048590422392
Gyc3_141 y3 0 x141 0 0.0201331642526096
Gyc3_142 y3 0 x142 0 -0.0515015627777372
Gyc3_143 y3 0 x143 0 0.0597284060510588
Gyc3_144 y3 0 x144 0 0.020165026634466
Gyc3_145 y3 0 x145 0 -0.0172858036775518
Gyc3_146 y3 0 x146 0 -0.0533354735065421
Gyc3_147 y3 0 x147 0 0.10048948561623
Gyc3_148 y3 0 x148 0 0.0720675991605814
Gyc3_149 y3 0 x149 0 -0.0240176249177025
Gyc3_150 y3 0 x150 0 -0.218177206623723
Gyc3_151 y3 0 x151 0 -0.0219137741534188
Gyc3_152 y3 0 x152 0 -0.0825993064349736
Gyc3_153 y3 0 x153 0 -0.0129133815767741
Gyc3_154 y3 0 x154 0 -0.00565313612722591
Gyc3_155 y3 0 x155 0 0.196107062145214
Gyc3_156 y3 0 x156 0 0.0120239910274266
Gyc3_157 y3 0 x157 0 0.18601505750784
Gyc3_158 y3 0 x158 0 0.076293596491273
Gyc3_159 y3 0 x159 0 -0.00501862954085573
Gyc3_160 y3 0 x160 0 0.0138399158737786
Gyc3_161 y3 0 x161 0 -0.0236954758769639
Gyc3_162 y3 0 x162 0 0.0019622503572326
Gyc3_163 y3 0 x163 0 0.0415710742652717
Gyc3_164 y3 0 x164 0 -0.113127741693978
Gyc3_165 y3 0 x165 0 -0.00793278499433122
Gyc3_166 y3 0 x166 0 0.0575009339470277
Gyc3_167 y3 0 x167 0 0.0703154515605427
Gyc3_168 y3 0 x168 0 0.0387929600724192
Gyc3_169 y3 0 x169 0 0.110550156437492
Gyc3_170 y3 0 x170 0 -0.0348394735714762
Gyc3_171 y3 0 x171 0 0.463761318323468
Gyc3_172 y3 0 x172 0 0.0725148786006533
Gyc3_173 y3 0 x173 0 -0.0314671833282738
Gyc3_174 y3 0 x174 0 0.0339079314210027
Gyc3_175 y3 0 x175 0 0.0816732398315501
Gyc3_176 y3 0 x176 0 -0.00729011296368055
Gyc3_177 y3 0 x177 0 -0.0825681490620722
Gyc3_178 y3 0 x178 0 -0.00497565974840429
Gyc3_179 y3 0 x179 0 0.25198400707866
Gyc3_180 y3 0 x180 0 0.0558787706097022
Gyc3_181 y3 0 x181 0 0.0943189406449485
Gyc3_182 y3 0 x182 0 0.0167114824387288
Gyc3_183 y3 0 x183 0 0.0394123374002712
Gyc3_184 y3 0 x184 0 -0.0394639041639914
Gyc3_185 y3 0 x185 0 -0.0036156873598767
Gyc3_186 y3 0 x186 0 -0.00967204628330308
Gyc3_187 y3 0 x187 0 -0.0216794418145788
Gyc3_188 y3 0 x188 0 -0.0264222208204208
Gyc3_189 y3 0 x189 0 0.0399568900710807
Gyc3_190 y3 0 x190 0 -0.118652755234882
Gyc3_191 y3 0 x191 0 -0.0378983353799671
Gyc3_192 y3 0 x192 0 0.105809774262424
Gyc3_193 y3 0 x193 0 -0.275516287175673
Gyc3_194 y3 0 x194 0 0.000140191857904571
Gyc3_195 y3 0 x195 0 0.0265867132886568
Gyc3_196 y3 0 x196 0 0.00330127500639541
Gyc3_197 y3 0 x197 0 -0.100469507682243
Gyc3_198 y3 0 x198 0 -0.187783247285866
Gyc3_199 y3 0 x199 0 -0.499302264601164
Gyc3_200 y3 0 x200 0 -0.487882808128295
Gyc3_201 y3 0 x201 0 -1
Gyc3_202 y3 0 x202 0 0.569157441024388
Gyc3_203 y3 0 x203 0 -0.502250944715357
Gyc3_204 y3 0 x204 0 0.927922460528624
Gyc3_205 y3 0 x205 0 -0.340844162277694
Gyc3_206 y3 0 x206 0 0.535610346967597
Gyc3_207 y3 0 x207 0 -0.90672147598372
Gyc3_208 y3 0 x208 0 0.0326132862866933
Gyc3_209 y3 0 x209 0 -0.241136824614316
Gyc3_210 y3 0 x210 0 -1
Gyc3_211 y3 0 x211 0 -0.887285852355571
Gyc3_212 y3 0 x212 0 -0.26067359768789
Gyc3_213 y3 0 x213 0 -0.33156876388218
Gyc3_214 y3 0 x214 0 -1
Gyc3_215 y3 0 x215 0 1
Gyc3_216 y3 0 x216 0 0.212682012119214
Gyc3_217 y3 0 x217 0 1
Gyc3_218 y3 0 x218 0 -0.644369559009898
Gyc3_219 y3 0 x219 0 0.795471772696244
Gyc3_220 y3 0 x220 0 -0.0342180309324703
Gyc3_221 y3 0 x221 0 0.136351926416886
Gyc3_222 y3 0 x222 0 1
Gyc3_223 y3 0 x223 0 0.0354280695030493
Gyc3_224 y3 0 x224 0 0.896546360897508
Gyc3_225 y3 0 x225 0 -0.095918302501703
Gyc3_226 y3 0 x226 0 1
Gyc3_227 y3 0 x227 0 0.839832251926193
Gyc3_228 y3 0 x228 0 -0.148670329553687
Gyc3_229 y3 0 x229 0 -1
Gyc3_230 y3 0 x230 0 -0.144126868139507
Gyc3_231 y3 0 x231 0 0.0679230940759598
Gyc3_232 y3 0 x232 0 -1
Gyc3_233 y3 0 x233 0 0.961247987674824
Gyc3_234 y3 0 x234 0 0.311761901740297
Gyc3_235 y3 0 x235 0 0.954307959380036
Gyc3_236 y3 0 x236 0 -0.790409580232169
Gyc3_237 y3 0 x237 0 -0.513562698304707
Gyc3_238 y3 0 x238 0 1
Gyc3_239 y3 0 x239 0 0.199849002379436
Gyc3_240 y3 0 x240 0 -0.925408264474808
Gyc3_241 y3 0 x241 0 0.879200802794141
Gyc3_242 y3 0 x242 0 0.0365624927768198
Gyc3_243 y3 0 x243 0 0.197513731461824
Gyc3_244 y3 0 x244 0 1
Gyc3_245 y3 0 x245 0 -0.0190601310364466
Gyc3_246 y3 0 x246 0 1
Gyc3_247 y3 0 x247 0 0.71021334071166
Gyc3_248 y3 0 x248 0 1
Gyc3_249 y3 0 x249 0 1
Gyc3_250 y3 0 x250 0 1
Gyc3_251 y3 0 x251 0 -0.548152338399761
Gyc3_252 y3 0 x252 0 0.56361922925226
Gyc3_253 y3 0 x253 0 -1
Gyc3_254 y3 0 x254 0 -0.496814934137457
Gyc3_255 y3 0 x255 0 -1
Gyc3_256 y3 0 x256 0 1
Gyc3_257 y3 0 x257 0 0.200116094454055
Gyc3_258 y3 0 x258 0 -1
Gyc3_259 y3 0 x259 0 -1
Gyc3_260 y3 0 x260 0 -0.672337292184254
Gyc3_261 y3 0 x261 0 0.242999608903781
Gyc3_262 y3 0 x262 0 0.37878833705752
Gyc3_263 y3 0 x263 0 -1
Gyc3_264 y3 0 x264 0 -1
Gyc3_265 y3 0 x265 0 0.0668339177713878
Gyc3_266 y3 0 x266 0 0.840495507234262
Gyc3_267 y3 0 x267 0 0.6680462797895
Gyc3_268 y3 0 x268 0 0.692935793122098
Gyc3_269 y3 0 x269 0 -1
Gyc3_270 y3 0 x270 0 0.766358139246178
Gyc3_271 y3 0 x271 0 -0.682681546806899
Gyc3_272 y3 0 x272 0 0.423762694010253
Gyc3_273 y3 0 x273 0 -0.930277425708249
Gyc3_274 y3 0 x274 0 -0.0450736777172147
Gyc3_275 y3 0 x275 0 -0.873220959423369
Gyc3_276 y3 0 x276 0 -1
Gyc3_277 y3 0 x277 0 0.539825057791194
Gyc3_278 y3 0 x278 0 -0.903530483196677
Gyc3_279 y3 0 x279 0 -1
Gyc3_280 y3 0 x280 0 -1
Gyc3_281 y3 0 x281 0 -0.0752312734843167
Gyc3_282 y3 0 x282 0 1
Gyc3_283 y3 0 x283 0 -1
Gyc3_284 y3 0 x284 0 0.617229600095199
Gyc3_285 y3 0 x285 0 -0.0906317932515045
Gyc3_286 y3 0 x286 0 -0.775905897925876
Gyc3_287 y3 0 x287 0 0.464909128001293
Gyc3_288 y3 0 x288 0 -0.953393758308521
Gyc3_289 y3 0 x289 0 1
Gyc3_290 y3 0 x290 0 -1
Gyc3_291 y3 0 x291 0 0.0622204589582379
Gyc3_292 y3 0 x292 0 -0.246334955096598
Gyc3_293 y3 0 x293 0 1
Gyc3_294 y3 0 x294 0 0.520062305746319
Gyc3_295 y3 0 x295 0 0.311700402331977
Gyc3_296 y3 0 x296 0 0.0233068588827313
Gyc3_297 y3 0 x297 0 -0.736246928327315
Gyc3_298 y3 0 x298 0 0.809735976495283
Gyc3_299 y3 0 x299 0 -1
Gyc3_300 y3 0 x300 0 0.12760280331758
Gyc3_301 y3 0 x301 0 -1
Gyc3_302 y3 0 x302 0 0.788616935353728
Gyc3_303 y3 0 x303 0 -1
Gyc3_304 y3 0 x304 0 0.898425570399979
Gyc3_305 y3 0 x305 0 -0.160869086938189
Gyc3_306 y3 0 x306 0 -0.19923909044824
Gyc3_307 y3 0 x307 0 -1
Gyc3_308 y3 0 x308 0 -0.284729275061268
Gyc3_309 y3 0 x309 0 1
Gyc3_310 y3 0 x310 0 -0.492672184155851
Gyc3_311 y3 0 x311 0 1
Gyc3_312 y3 0 x312 0 -0.333629317184589
Gyc3_313 y3 0 x313 0 1
Gyc3_314 y3 0 x314 0 1
Gyc3_315 y3 0 x315 0 -0.289638576563341
Gyc3_316 y3 0 x316 0 -0.158174810771842
Gyc3_317 y3 0 x317 0 0.21748382395963
Gyc3_318 y3 0 x318 0 0.68401876853848
Gyc3_319 y3 0 x319 0 0.842429935969754
Gyc3_320 y3 0 x320 0 -1
Gyc3_321 y3 0 x321 0 1
Gyc3_322 y3 0 x322 0 0.852513343007846
Gyc3_323 y3 0 x323 0 1
Gyc3_324 y3 0 x324 0 1
Gyc3_325 y3 0 x325 0 1
Gyc3_326 y3 0 x326 0 -1
Gyc3_327 y3 0 x327 0 -0.501812507241219
Gyc3_328 y3 0 x328 0 -0.648550790951506
Gyc3_329 y3 0 x329 0 -1
Gyc3_330 y3 0 x330 0 0.416777310686901
Gyc3_331 y3 0 x331 0 -1
Gyc3_332 y3 0 x332 0 -1
Gyc3_333 y3 0 x333 0 0.801891025913485
Gyc3_334 y3 0 x334 0 1
Gyc3_335 y3 0 x335 0 0.206688450218613
Gyc3_336 y3 0 x336 0 0.419489795619584
Gyc3_337 y3 0 x337 0 1
Gyc3_338 y3 0 x338 0 -1
Gyc3_339 y3 0 x339 0 0.529690268616753
Gyc3_340 y3 0 x340 0 -1
Gyc3_341 y3 0 x341 0 1
Gyc3_342 y3 0 x342 0 -1
Gyc3_343 y3 0 x343 0 0.91067664973472
Gyc3_344 y3 0 x344 0 1
Gyc3_345 y3 0 x345 0 -0.165241100190688
Gyc3_346 y3 0 x346 0 -1
Gyc3_347 y3 0 x347 0 0.265082515746638
Gyc3_348 y3 0 x348 0 0.690790208541535
Gyc3_349 y3 0 x349 0 -1
Gyc3_350 y3 0 x350 0 -0.828239243928735
Gyc3_351 y3 0 x351 0 -1
Gyc3_352 y3 0 x352 0 0.304462495819207
Gyc3_353 y3 0 x353 0 -1
Gyc3_354 y3 0 x354 0 0.0638513583558362
Gyc3_355 y3 0 x355 0 0.340851546601434
Gyc3_356 y3 0 x356 0 -1
Gyc3_357 y3 0 x357 0 -0.130783356128206
Gyc3_358 y3 0 x358 0 1
Gyc3_359 y3 0 x359 0 -1
Gyc3_360 y3 0 x360 0 1
Gyc3_361 y3 0 x361 0 -1
Gyc3_362 y3 0 x362 0 -1
Gyc3_363 y3 0 x363 0 1
Gyc3_364 y3 0 x364 0 -1
Gyc3_365 y3 0 x365 0 0.976534238385832
Gyc3_366 y3 0 x366 0 1
Gyc3_367 y3 0 x367 0 0.640423174325508
Gyc3_368 y3 0 x368 0 1
Gyc3_369 y3 0 x369 0 -0.00189035655152874
Gyc3_370 y3 0 x370 0 -1
Gyc3_371 y3 0 x371 0 -0.0182843270687401
Gyc3_372 y3 0 x372 0 1
Gyc3_373 y3 0 x373 0 -1
Gyc3_374 y3 0 x374 0 1
Gyc3_375 y3 0 x375 0 1
Gyc3_376 y3 0 x376 0 -1
Gyc3_377 y3 0 x377 0 -1
Gyc3_378 y3 0 x378 0 -1
Gyc3_379 y3 0 x379 0 -0.595053077622719
Gyc3_380 y3 0 x380 0 1
Gyc3_381 y3 0 x381 0 1
Gyc3_382 y3 0 x382 0 1
Gyc3_383 y3 0 x383 0 1
Gyc3_384 y3 0 x384 0 -1
Gyc3_385 y3 0 x385 0 -1
Gyc3_386 y3 0 x386 0 -1
Gyc3_387 y3 0 x387 0 -0.912436118626062
Gyc3_388 y3 0 x388 0 -1
Gyc3_389 y3 0 x389 0 1
Gyc3_390 y3 0 x390 0 -0.492810174096319
Gyc3_391 y3 0 x391 0 -1
Gyc3_392 y3 0 x392 0 0.829627956838195
Gyc3_393 y3 0 x393 0 -1
Gyc3_394 y3 0 x394 0 -1
Gyc3_395 y3 0 x395 0 0.0283048688499825
Gyc3_396 y3 0 x396 0 1
Gyc3_397 y3 0 x397 0 1
Gyc3_398 y3 0 x398 0 -0.264460863658181
Gyc3_399 y3 0 x399 0 0.517358141776322
Gyc3_400 y3 0 x400 0 0.701640036894701
Gyc3_401 y3 0 x401 0 -1
Gyc3_402 y3 0 x402 0 1
Gyc3_403 y3 0 x403 0 1
Gyc3_404 y3 0 x404 0 1
Gyc3_405 y3 0 x405 0 1
Gyc3_406 y3 0 x406 0 1
Gyc3_407 y3 0 x407 0 -0.538078518420002
Gyc3_408 y3 0 x408 0 1
Gyc3_409 y3 0 x409 0 -1
Gyc3_410 y3 0 x410 0 1
Gyc3_411 y3 0 x411 0 -1
Gyc3_412 y3 0 x412 0 1
Gyc3_413 y3 0 x413 0 -1
Gyc3_414 y3 0 x414 0 -1
Gyc3_415 y3 0 x415 0 -1
Gyc3_416 y3 0 x416 0 -1
Gyc3_417 y3 0 x417 0 -1
Gyc3_418 y3 0 x418 0 -1
Gyc3_419 y3 0 x419 0 1
Gyc3_420 y3 0 x420 0 -1
Gyc3_421 y3 0 x421 0 1
Gyc3_422 y3 0 x422 0 -1
Gyc3_423 y3 0 x423 0 1
Gyc3_424 y3 0 x424 0 1
Gyc3_425 y3 0 x425 0 1
Gyc3_426 y3 0 x426 0 1
Gyc3_427 y3 0 x427 0 1
Gyc3_428 y3 0 x428 0 -1
Gyc3_429 y3 0 x429 0 -1
Gyc3_430 y3 0 x430 0 1
Gyc3_431 y3 0 x431 0 -1
Gyc3_432 y3 0 x432 0 -1
Gyc3_433 y3 0 x433 0 1
Gyc3_434 y3 0 x434 0 -1
Gyc3_435 y3 0 x435 0 -1
Gyc3_436 y3 0 x436 0 -1
Gyc3_437 y3 0 x437 0 1
Gyc3_438 y3 0 x438 0 1
Gyc3_439 y3 0 x439 0 -1
Gyc3_440 y3 0 x440 0 -1
Gyc3_441 y3 0 x441 0 1
Gyc3_442 y3 0 x442 0 -1
Gyc3_443 y3 0 x443 0 1
Gyc3_444 y3 0 x444 0 1
Gyc3_445 y3 0 x445 0 1
Gyc3_446 y3 0 x446 0 1
Gyc3_447 y3 0 x447 0 1
Gyc3_448 y3 0 x448 0 -1
Gyc3_449 y3 0 x449 0 1
Gyc3_450 y3 0 x450 0 1
Gyc3_451 y3 0 x451 0 0.450149248638242
Gyc3_452 y3 0 x452 0 1
Gyc3_453 y3 0 x453 0 -1
Gyc3_454 y3 0 x454 0 1
Gyc3_455 y3 0 x455 0 0.686217874084557
Gyc3_456 y3 0 x456 0 1
Gyc3_457 y3 0 x457 0 -1
Gyc3_458 y3 0 x458 0 -1
Gyc3_459 y3 0 x459 0 -1
Gyc3_460 y3 0 x460 0 0.883288861910785
Gyc3_461 y3 0 x461 0 1
Gyc3_462 y3 0 x462 0 -1
Gyc3_463 y3 0 x463 0 -1
Gyc3_464 y3 0 x464 0 0.749228753521753
Gyc3_465 y3 0 x465 0 1
Gyc3_466 y3 0 x466 0 1
Gyc3_467 y3 0 x467 0 1
Gyc3_468 y3 0 x468 0 1
Gyc3_469 y3 0 x469 0 -1
Gyc3_470 y3 0 x470 0 1
Gyc3_471 y3 0 x471 0 -0.484301624234549
Gyc3_472 y3 0 x472 0 1
Gyc3_473 y3 0 x473 0 -1
Gyc3_474 y3 0 x474 0 0.305129536138071
Gyc3_475 y3 0 x475 0 -1
Gyc3_476 y3 0 x476 0 1
Gyc3_477 y3 0 x477 0 1
Gyc3_478 y3 0 x478 0 -1
Gyc3_479 y3 0 x479 0 -1
Gyc3_480 y3 0 x480 0 -1
Gyc3_481 y3 0 x481 0 1
Gyc3_482 y3 0 x482 0 1
Gyc3_483 y3 0 x483 0 -1
Gyc3_484 y3 0 x484 0 0.61877239903927
Gyc3_485 y3 0 x485 0 -1
Gyc3_486 y3 0 x486 0 -1
Gyc3_487 y3 0 x487 0 1
Gyc3_488 y3 0 x488 0 -1
Gyc3_489 y3 0 x489 0 1
Gyc3_490 y3 0 x490 0 -1
Gyc3_491 y3 0 x491 0 1
Gyc3_492 y3 0 x492 0 -1
Gyc3_493 y3 0 x493 0 1
Gyc3_494 y3 0 x494 0 -0.0143220430203132
Gyc3_495 y3 0 x495 0 1
Gyc3_496 y3 0 x496 0 1
Gyc3_497 y3 0 x497 0 1
Gyc3_498 y3 0 x498 0 1
Gyc3_499 y3 0 x499 0 1
Gyc3_500 y3 0 x500 0 1
Gyc3_501 y3 0 x501 0 -0.488447575770873
Gyc3_502 y3 0 x502 0 1
Gyc3_503 y3 0 x503 0 -0.082036972638291
Gyc3_504 y3 0 x504 0 1
Gyc3_505 y3 0 x505 0 1
Gyc3_506 y3 0 x506 0 -1
Gyc3_507 y3 0 x507 0 -1
Gyc3_508 y3 0 x508 0 1
Gyc3_509 y3 0 x509 0 0.637209085955649
Gyc3_510 y3 0 x510 0 -1
Gyc3_511 y3 0 x511 0 1
Gyc3_512 y3 0 x512 0 -1
Gyc3_513 y3 0 x513 0 1
Gyc3_514 y3 0 x514 0 1
Gyc3_515 y3 0 x515 0 -1
Gyc3_516 y3 0 x516 0 1
Gyc3_517 y3 0 x517 0 1
Gyc3_518 y3 0 x518 0 1
Gyc3_519 y3 0 x519 0 -1
Gyc3_520 y3 0 x520 0 1
Gyc3_521 y3 0 x521 0 1
Gyc3_522 y3 0 x522 0 1
Gyc3_523 y3 0 x523 0 0.314943157193031
Gyc3_524 y3 0 x524 0 1
Gyc3_525 y3 0 x525 0 1
Gyc3_526 y3 0 x526 0 -1
Gyc3_527 y3 0 x527 0 1
Gyc3_528 y3 0 x528 0 -1
Gyc3_529 y3 0 x529 0 -1
Gyc3_530 y3 0 x530 0 -1
Gyc3_531 y3 0 x531 0 -1
Gyc3_532 y3 0 x532 0 -1
Gyc3_533 y3 0 x533 0 1
Gyc3_534 y3 0 x534 0 1
Gyc3_535 y3 0 x535 0 -1
Gyc3_536 y3 0 x536 0 1
Gyc3_537 y3 0 x537 0 1
Gyc3_538 y3 0 x538 0 -1
Gyc3_539 y3 0 x539 0 1
Gyc3_540 y3 0 x540 0 0.746365002306818
Gyc3_541 y3 0 x541 0 1
Gyc3_542 y3 0 x542 0 -1
Gyc3_543 y3 0 x543 0 1
Gyc3_544 y3 0 x544 0 1
Gyc3_545 y3 0 x545 0 -1
Gyc3_546 y3 0 x546 0 -1
Gyc3_547 y3 0 x547 0 1
Gyc3_548 y3 0 x548 0 -1
Gyc3_549 y3 0 x549 0 -1
Gyc3_550 y3 0 x550 0 -1
Gyc3_551 y3 0 x551 0 -1
Gyc3_552 y3 0 x552 0 -1
Gyc3_553 y3 0 x553 0 -1
Gyc3_554 y3 0 x554 0 -1
Gyc3_555 y3 0 x555 0 -1
Gyc3_556 y3 0 x556 0 -1
Gyc3_557 y3 0 x557 0 1
Gyc3_558 y3 0 x558 0 0.648977195181731
Gyc3_559 y3 0 x559 0 -1
Gyc3_560 y3 0 x560 0 -0.465470806707079
Gyc3_561 y3 0 x561 0 -1
Gyc3_562 y3 0 x562 0 -1
Gyc3_563 y3 0 x563 0 1
Gyc3_564 y3 0 x564 0 -1
Gyc3_565 y3 0 x565 0 1
Gyc3_566 y3 0 x566 0 1
Gyc3_567 y3 0 x567 0 1
Gyc3_568 y3 0 x568 0 1
Gyc3_569 y3 0 x569 0 -1
Gyc3_570 y3 0 x570 0 -1
Gyc3_571 y3 0 x571 0 1
Gyc3_572 y3 0 x572 0 1
Gyc3_573 y3 0 x573 0 -1
Gyc3_574 y3 0 x574 0 1
Gyc3_575 y3 0 x575 0 -1
Gyc3_576 y3 0 x576 0 -1
Gyc3_577 y3 0 x577 0 -1
Gyc3_578 y3 0 x578 0 -1
Gyc3_579 y3 0 x579 0 1
Gyc3_580 y3 0 x580 0 1
Gyc3_581 y3 0 x581 0 1
Gyc3_582 y3 0 x582 0 1
Gyc3_583 y3 0 x583 0 1
Gyc3_584 y3 0 x584 0 -1
Gyc3_585 y3 0 x585 0 -1
Gyc3_586 y3 0 x586 0 -0.220140981431934
Gyc3_587 y3 0 x587 0 -1
Gyc3_588 y3 0 x588 0 -1
Gyc3_589 y3 0 x589 0 1
Gyc3_590 y3 0 x590 0 -1
Gyc3_591 y3 0 x591 0 -1
Gyc3_592 y3 0 x592 0 1
Gyc3_593 y3 0 x593 0 -1
Gyc3_594 y3 0 x594 0 -1
Gyc3_595 y3 0 x595 0 1
Gyc3_596 y3 0 x596 0 1
Gyc3_597 y3 0 x597 0 0.161769881990142
Gyc3_598 y3 0 x598 0 -1
Gyc3_599 y3 0 x599 0 1
Gyc3_600 y3 0 x600 0 1
Gyd3_1 y3 0 u1 0 -0.276371351645904
Gyd3_2 y3 0 u2 0 -0.568346326707177
Gyd3_3 y3 0 u3 0 -3.6536002292946
.ENDS
