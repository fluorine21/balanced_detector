* Equivalent circuit model for HMC539ALP3E_4dB.ckt
.SUBCKT HMC539ALP3E_4dB po1 po2
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Vsp2 po2 p2 0
Vsr2 p2 pr2 0
Rp2 pr2 0 50
Ru2 u2 0 50
Fr2 u2 0 Vsr2 -1
Fu2 u2 0 Vsp2 -1
Ry2 y2 0 1
Gy2 p2 0 y2 0 -0.02
Rx1 x1 0 1
Cx1 x1 0 3.53627063161835e-13
Gx1_1 x1 0 u1 0 -23.3354738307188
Rx2 x2 0 1
Cx2 x2 0 8.59855014759414e-12
Gx2_1 x2 0 u1 0 -146.195139162122
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 96.5889608593002
Cx3 x3 xm3 1.52013265599724e-13
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -0.0143272903577363
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -84.6791663726074
Cx4 x4 xm4 1.52013265599724e-13
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 1.2132230038714
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 19.7968365880108
Cx5 x5 xm5 1.34030288980988e-11
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -123.828239960321
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -0.0298487059512434
Cx6 x6 xm6 1.34030288980988e-11
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 3.69611272303563
Rx7 x7 0 1
Fxc7_8 x7 0 Vx8 303.516760110041
Cx7 x7 xm7 3.10934658884836e-14
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 -2.32735882357128e-07
Rx8 x8 0 1
Fxc8_7 x8 0 Vx7 -866.471687313706
Cx8 x8 xm8 3.10934658884836e-14
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 0.000201659052684425
Rx9 x9 0 1
Fxc9_10 x9 0 Vx10 7621.61474146488
Cx9 x9 xm9 8.40733664871429e-15
Vx9 xm9 0 0
Gx9_1 x9 0 u1 0 -1.60216415289659e-08
Rx10 x10 0 1
Fxc10_9 x10 0 Vx9 -476.66364935604
Cx10 x10 xm10 8.40733664871429e-15
Vx10 xm10 0 0
Gx10_1 x10 0 u1 0 7.63693411987119e-06
Rx11 x11 0 1
Fxc11_12 x11 0 Vx12 31466.3025109729
Cx11 x11 xm11 1.94523784543502e-15
Vx11 xm11 0 0
Gx11_1 x11 0 u1 0 -3.14096139534946e-10
Rx12 x12 0 1
Fxc12_11 x12 0 Vx11 -2166.3912177589
Cx12 x12 xm12 1.94523784543502e-15
Vx12 xm12 0 0
Gx12_1 x12 0 u1 0 6.80455118220479e-07
Rx13 x13 0 1
Fxc13_14 x13 0 Vx14 276.511576551915
Cx13 x13 xm13 1.91730724654873e-14
Vx13 xm13 0 0
Gx13_1 x13 0 u1 0 -2.64181685207841e-08
Rx14 x14 0 1
Fxc14_13 x14 0 Vx13 -2554.77379077861
Cx14 x14 xm14 1.91730724654873e-14
Vx14 xm14 0 0
Gx14_1 x14 0 u1 0 6.7492444537272e-05
Rx15 x15 0 1
Fxc15_16 x15 0 Vx16 138.773612037799
Cx15 x15 xm15 4.56584091846018e-14
Vx15 xm15 0 0
Gx15_1 x15 0 u1 0 -3.01357776271498e-07
Rx16 x16 0 1
Fxc16_15 x16 0 Vx15 -903.198020640163
Cx16 x16 xm16 4.56584091846018e-14
Vx16 xm16 0 0
Gx16_1 x16 0 u1 0 0.000272185747032938
Rx17 x17 0 1
Fxc17_18 x17 0 Vx18 124666.448398836
Cx17 x17 xm17 6.22970485029519e-16
Vx17 xm17 0 0
Gx17_1 x17 0 u1 0 -1.81171897085339e-10
Rx18 x18 0 1
Fxc18_17 x18 0 Vx17 -5426.52487040467
Cx18 x18 xm18 6.22970485029519e-16
Vx18 xm18 0 0
Gx18_1 x18 0 u1 0 9.83133805351986e-07
Rx19 x19 0 1
Fxc19_20 x19 0 Vx20 17.5112589039375
Cx19 x19 xm19 1.1019165711965e-12
Vx19 xm19 0 0
Gx19_1 x19 0 u1 0 -0.0616832679103059
Rx20 x20 0 1
Fxc20_19 x20 0 Vx19 -13.6596549192874
Cx20 x20 xm20 1.1019165711965e-12
Vx20 xm20 0 0
Gx20_1 x20 0 u1 0 0.842572153948733
Rx21 x21 0 1
Fxc21_22 x21 0 Vx22 41923.3982965501
Cx21 x21 xm21 4.28178588649374e-16
Vx21 xm21 0 0
Gx21_1 x21 0 u1 0 -2.11246259241297e-10
Rx22 x22 0 1
Fxc22_21 x22 0 Vx21 -34421.1379400114
Cx22 x22 xm22 4.28178588649374e-16
Vx22 xm22 0 0
Gx22_1 x22 0 u1 0 7.27133662865608e-06
Rx23 x23 0 1
Fxc23_24 x23 0 Vx24 3611.81981174937
Cx23 x23 xm23 2.43387977270851e-14
Vx23 xm23 0 0
Gx23_1 x23 0 u1 0 -1.27205224656701e-07
Rx24 x24 0 1
Fxc24_23 x24 0 Vx23 -124.040656070295
Cx24 x24 xm24 2.43387977270851e-14
Vx24 xm24 0 0
Gx24_1 x24 0 u1 0 1.57786195219864e-05
Rx25 x25 0 1
Fxc25_26 x25 0 Vx26 101.367453795337
Cx25 x25 xm25 1.05011663800036e-13
Vx25 xm25 0 0
Gx25_1 x25 0 u1 0 -5.90736051735668e-06
Rx26 x26 0 1
Fxc26_25 x26 0 Vx25 -239.324004079753
Cx26 x26 xm26 1.05011663800036e-13
Vx26 xm26 0 0
Gx26_1 x26 0 u1 0 0.00141377317255644
Rx27 x27 0 1
Fxc27_28 x27 0 Vx28 132.701314661351
Cx27 x27 xm27 1.08883637079586e-14
Vx27 xm27 0 0
Gx27_1 x27 0 u1 0 -1.46671824042291e-09
Rx28 x28 0 1
Fxc28_27 x28 0 Vx27 -17125.4555074516
Cx28 x28 xm28 1.08883637079586e-14
Vx28 xm28 0 0
Gx28_1 x28 0 u1 0 2.51182179683303e-05
Rx29 x29 0 1
Fxc29_30 x29 0 Vx30 686.732174778935
Cx29 x29 xm29 1.79569174984714e-14
Vx29 xm29 0 0
Gx29_1 x29 0 u1 0 -4.02991480661098e-08
Rx30 x30 0 1
Fxc30_29 x30 0 Vx29 -1223.40114623618
Cx30 x30 xm30 1.79569174984714e-14
Vx30 xm30 0 0
Gx30_1 x30 0 u1 0 4.930202393642e-05
Rx31 x31 0 1
Fxc31_32 x31 0 Vx32 705.853631531373
Cx31 x31 xm31 1.89102617067545e-14
Vx31 xm31 0 0
Gx31_1 x31 0 u1 0 -4.48220061496545e-08
Rx32 x32 0 1
Fxc32_31 x32 0 Vx31 -1078.69458135216
Cx32 x32 xm32 1.89102617067545e-14
Vx32 xm32 0 0
Gx32_1 x32 0 u1 0 4.83492551589656e-05
Rx33 x33 0 1
Fxc33_34 x33 0 Vx34 3398.42629107471
Cx33 x33 xm33 1.08306461059872e-14
Vx33 xm33 0 0
Gx33_1 x33 0 u1 0 -1.44661884383519e-08
Rx34 x34 0 1
Fxc34_33 x34 0 Vx33 -686.794643951847
Cx34 x34 xm34 1.08306461059872e-14
Vx34 xm34 0 0
Gx34_1 x34 0 u1 0 9.93530073785823e-06
Rx35 x35 0 1
Fxc35_36 x35 0 Vx36 32.9195435907089
Cx35 x35 xm35 2.09659001892218e-13
Vx35 xm35 0 0
Gx35_1 x35 0 u1 0 -0.000130411267904078
Rx36 x36 0 1
Fxc36_35 x36 0 Vx35 -193.726420201423
Cx36 x36 xm36 2.09659001892218e-13
Vx36 xm36 0 0
Gx36_1 x36 0 u1 0 0.0252641080849858
Rx37 x37 0 1
Fxc37_38 x37 0 Vx38 1682.96727439499
Cx37 x37 xm37 1.6602740464064e-14
Vx37 xm37 0 0
Gx37_1 x37 0 u1 0 -2.47485809847296e-08
Rx38 x38 0 1
Fxc38_37 x38 0 Vx37 -597.485703431046
Cx38 x38 xm38 1.6602740464064e-14
Vx38 xm38 0 0
Gx38_1 x38 0 u1 0 1.47869233185814e-05
Rx39 x39 0 1
Fxc39_40 x39 0 Vx40 476.164953784541
Cx39 x39 xm39 1.17924667928284e-12
Vx39 xm39 0 0
Gx39_1 x39 0 u1 0 -0.189260043541653
Rx40 x40 0 1
Fxc40_39 x40 0 Vx39 -0.489820742772458
Cx40 x40 xm40 1.17924667928284e-12
Vx40 xm40 0 0
Gx40_1 x40 0 u1 0 0.0927034951047201
Rx41 x41 0 1
Fxc41_42 x41 0 Vx42 47.2049658983037
Cx41 x41 xm41 2.25551329603533e-13
Vx41 xm41 0 0
Gx41_1 x41 0 u1 0 -0.000242737201493873
Rx42 x42 0 1
Fxc42_41 x42 0 Vx41 -117.762215125279
Cx42 x42 xm42 2.25551329603533e-13
Vx42 xm42 0 0
Gx42_1 x42 0 u1 0 0.0285852705412296
Rx43 x43 0 1
Fxc43_44 x43 0 Vx44 2217.78939647574
Cx43 x43 xm43 3.84602500012975e-15
Vx43 xm43 0 0
Gx43_1 x43 0 u1 0 -1.01835111571991e-09
Rx44 x44 0 1
Fxc44_43 x44 0 Vx43 -8495.42422056443
Cx44 x44 xm44 3.84602500012975e-15
Vx44 xm44 0 0
Gx44_1 x44 0 u1 0 8.65132473352573e-06
Rx45 x45 0 1
Fxc45_46 x45 0 Vx46 5797.91647742002
Cx45 x45 xm45 9.27706506013979e-15
Vx45 xm45 0 0
Gx45_1 x45 0 u1 0 -9.45866302498017e-09
Rx46 x46 0 1
Fxc46_45 x46 0 Vx45 -563.577085646458
Cx46 x46 xm46 9.27706506013979e-15
Vx46 xm46 0 0
Gx46_1 x46 0 u1 0 5.33068574173024e-06
Rx47 x47 0 1
Fxc47_48 x47 0 Vx48 9871.13909251475
Cx47 x47 xm47 2.25851726135813e-15
Vx47 xm47 0 0
Gx47_1 x47 0 u1 0 -1.09585437116584e-09
Rx48 x48 0 1
Fxc48_47 x48 0 Vx47 -5629.32030229767
Cx48 x48 xm48 2.25851726135813e-15
Vx48 xm48 0 0
Gx48_1 x48 0 u1 0 6.16891525996549e-06
Rx49 x49 0 1
Fxc49_50 x49 0 Vx50 599.401121355322
Cx49 x49 xm49 3.37035623112366e-15
Vx49 xm49 0 0
Gx49_1 x49 0 u1 0 -3.32337891232732e-10
Rx50 x50 0 1
Fxc50_49 x50 0 Vx49 -42021.6872622546
Cx50 x50 xm50 3.37035623112366e-15
Vx50 xm50 0 0
Gx50_1 x50 0 u1 0 1.39653989307791e-05
Rx51 x51 0 1
Fxc51_52 x51 0 Vx52 553.124137716997
Cx51 x51 xm51 1.88174133254326e-14
Vx51 xm51 0 0
Gx51_1 x51 0 u1 0 -2.58257075907216e-08
Rx52 x52 0 1
Fxc52_51 x52 0 Vx51 -1466.44427570381
Cx52 x52 xm52 1.88174133254326e-14
Vx52 xm52 0 0
Gx52_1 x52 0 u1 0 3.78719610624142e-05
Rx53 x53 0 1
Fxc53_54 x53 0 Vx54 744.139564932269
Cx53 x53 xm53 1.207285936914e-14
Vx53 xm53 0 0
Gx53_1 x53 0 u1 0 -6.69318298580556e-09
Rx54 x54 0 1
Fxc54_53 x54 0 Vx53 -2666.66408656669
Cx54 x54 xm54 1.207285936914e-14
Vx54 xm54 0 0
Gx54_1 x54 0 u1 0 1.78484706930669e-05
Rx55 x55 0 1
Fxc55_56 x55 0 Vx56 3296.72413306488
Cx55 x55 xm55 1.59455172364102e-14
Vx55 xm55 0 0
Gx55_1 x55 0 u1 0 -1.38536433290349e-07
Rx56 x56 0 1
Fxc56_55 x56 0 Vx55 -348.125345022652
Cx56 x56 xm56 1.59455172364102e-14
Vx56 xm56 0 0
Gx56_1 x56 0 u1 0 4.82280436374105e-05
Rx57 x57 0 1
Fxc57_58 x57 0 Vx58 1444.7258862366
Cx57 x57 xm57 1.4256037936421e-14
Vx57 xm57 0 0
Gx57_1 x57 0 u1 0 -7.92138180885543e-08
Rx58 x58 0 1
Fxc58_57 x58 0 Vx57 -993.343810214827
Cx58 x58 xm58 1.4256037936421e-14
Vx58 xm58 0 0
Gx58_1 x58 0 u1 0 7.86865558817488e-05
Rx59 x59 0 1
Fxc59_60 x59 0 Vx60 91.7841654908644
Cx59 x59 xm59 1.54588556473979e-13
Vx59 xm59 0 0
Gx59_1 x59 0 u1 0 -1.7704566765159e-05
Rx60 x60 0 1
Fxc60_59 x60 0 Vx59 -135.366540724299
Cx60 x60 xm60 1.54588556473979e-13
Vx60 xm60 0 0
Gx60_1 x60 0 u1 0 0.00239660595802197
Rx61 x61 0 1
Fxc61_62 x61 0 Vx62 1175.9789421607
Cx61 x61 xm61 1.36270438718843e-15
Vx61 xm61 0 0
Gx61_1 x61 0 u1 0 -1.15562283929119e-11
Rx62 x62 0 1
Fxc62_61 x62 0 Vx61 -135174.510908694
Cx62 x62 xm62 1.36270438718843e-15
Vx62 xm62 0 0
Gx62_1 x62 0 u1 0 1.56210752096102e-06
Rx63 x63 0 1
Fxc63_64 x63 0 Vx64 275.384762980406
Cx63 x63 xm63 1.8842536609155e-14
Vx63 xm63 0 0
Gx63_1 x63 0 u1 0 -1.04777195177397e-08
Rx64 x64 0 1
Fxc64_63 x64 0 Vx63 -3032.8475700867
Cx64 x64 xm64 1.8842536609155e-14
Vx64 xm64 0 0
Gx64_1 x64 0 u1 0 3.17773261794268e-05
Rx65 x65 0 1
Fxc65_66 x65 0 Vx66 248.237264038468
Cx65 x65 xm65 2.58532363902921e-14
Vx65 xm65 0 0
Gx65_1 x65 0 u1 0 -3.37615437603464e-08
Rx66 x66 0 1
Fxc66_65 x66 0 Vx65 -1796.25712173453
Cx66 x66 xm66 2.58532363902921e-14
Vx66 xm66 0 0
Gx66_1 x66 0 u1 0 6.06444134202744e-05
Rx67 x67 0 1
Fxc67_68 x67 0 Vx68 6512.74600592457
Cx67 x67 xm67 4.40227995829476e-15
Vx67 xm67 0 0
Gx67_1 x67 0 u1 0 -1.4854945859221e-09
Rx68 x68 0 1
Fxc68_67 x68 0 Vx67 -2376.37011567801
Cx68 x68 xm68 4.40227995829476e-15
Vx68 xm68 0 0
Gx68_1 x68 0 u1 0 3.53008494098676e-06
Rx69 x69 0 1
Fxc69_70 x69 0 Vx70 1195.14057961071
Cx69 x69 xm69 2.0912663085398e-14
Vx69 xm69 0 0
Gx69_1 x69 0 u1 0 -4.11924789406929e-08
Rx70 x70 0 1
Fxc70_69 x70 0 Vx69 -578.551412630745
Cx70 x70 xm70 2.0912663085398e-14
Vx70 xm70 0 0
Gx70_1 x70 0 u1 0 2.38319668809001e-05
Rx71 x71 0 1
Fxc71_72 x71 0 Vx72 1082.09640680966
Cx71 x71 xm71 6.45713973054353e-15
Vx71 xm71 0 0
Gx71_1 x71 0 u1 0 -1.14044157455275e-09
Rx72 x72 0 1
Fxc72_71 x72 0 Vx71 -6758.38775284539
Cx72 x72 xm72 6.45713973054353e-15
Vx72 xm72 0 0
Gx72_1 x72 0 u1 0 7.707546370293e-06
Rx73 x73 0 1
Fxc73_74 x73 0 Vx74 1206.12578085641
Cx73 x73 xm73 7.88540425403586e-15
Vx73 xm73 0 0
Gx73_1 x73 0 u1 0 -1.15559666205946e-09
Rx74 x74 0 1
Fxc74_73 x74 0 Vx73 -4088.78232534124
Cx74 x74 xm74 7.88540425403586e-15
Vx74 xm74 0 0
Gx74_1 x74 0 u1 0 4.72498320705204e-06
Rx75 x75 0 1
Fxc75_76 x75 0 Vx76 61.6537369217556
Cx75 x75 xm75 1.62084283086177e-13
Vx75 xm75 0 0
Gx75_1 x75 0 u1 0 -1.01303717079158e-05
Rx76 x76 0 1
Fxc76_75 x76 0 Vx75 -201.70635215655
Cx76 x76 xm76 1.62084283086177e-13
Vx76 xm76 0 0
Gx76_1 x76 0 u1 0 0.00204336032319362
Rx77 x77 0 1
Fxc77_78 x77 0 Vx78 1686.83077689263
Cx77 x77 xm77 5.31549963067726e-14
Vx77 xm77 0 0
Gx77_1 x77 0 u1 0 -3.85153608469495e-07
Rx78 x78 0 1
Fxc78_77 x78 0 Vx77 -65.1882136985263
Cx78 x78 xm78 5.31549963067726e-14
Vx78 xm78 0 0
Gx78_1 x78 0 u1 0 2.5107475735668e-05
Rx79 x79 0 1
Fxc79_80 x79 0 Vx80 95.629611751479
Cx79 x79 xm79 1.78816112180161e-14
Vx79 xm79 0 0
Gx79_1 x79 0 u1 0 -2.23754529116245e-09
Rx80 x80 0 1
Fxc80_79 x80 0 Vx79 -10120.1990918297
Cx80 x80 xm80 1.78816112180161e-14
Vx80 xm80 0 0
Gx80_1 x80 0 u1 0 2.26444038235499e-05
Rx81 x81 0 1
Fxc81_82 x81 0 Vx82 1535.76946999461
Cx81 x81 xm81 7.76754927887759e-15
Vx81 xm81 0 0
Gx81_1 x81 0 u1 0 -3.38084315624999e-10
Rx82 x82 0 1
Fxc82_81 x82 0 Vx81 -3372.5035410279
Cx82 x82 xm82 7.76754927887759e-15
Vx82 xm82 0 0
Gx82_1 x82 0 u1 0 1.1401905516113e-06
Rx83 x83 0 1
Fxc83_84 x83 0 Vx84 21025.0722219935
Cx83 x83 xm83 1.25557410678191e-15
Vx83 xm83 0 0
Gx83_1 x83 0 u1 0 -6.68887450808163e-11
Rx84 x84 0 1
Fxc84_83 x84 0 Vx83 -9486.03810211623
Cx84 x84 xm84 1.25557410678191e-15
Vx84 xm84 0 0
Gx84_1 x84 0 u1 0 6.34509184439363e-07
Rx85 x85 0 1
Fxc85_86 x85 0 Vx86 681.323069053088
Cx85 x85 xm85 1.63787697489454e-14
Vx85 xm85 0 0
Gx85_1 x85 0 u1 0 -7.82250989938739e-09
Rx86 x86 0 1
Fxc86_85 x86 0 Vx85 -1789.60005859728
Cx86 x86 xm86 1.63787697489454e-14
Vx86 xm86 0 0
Gx86_1 x86 0 u1 0 1.39991641743215e-05
Rx87 x87 0 1
Fxc87_88 x87 0 Vx88 1708.08094626546
Cx87 x87 xm87 1.19981261746115e-15
Vx87 xm87 0 0
Gx87_1 x87 0 u1 0 -3.10458603563905e-11
Rx88 x88 0 1
Fxc88_87 x88 0 Vx87 -128626.540410533
Cx88 x88 xm88 1.19981261746115e-15
Vx88 xm88 0 0
Gx88_1 x88 0 u1 0 3.99332161171104e-06
Rx89 x89 0 1
Fxc89_90 x89 0 Vx90 286644.320976722
Cx89 x89 xm89 6.90011418477151e-16
Vx89 xm89 0 0
Gx89_1 x89 0 u1 0 -4.82826706878645e-10
Rx90 x90 0 1
Fxc90_89 x90 0 Vx89 -2385.8102256165
Cx90 x90 xm90 6.90011418477151e-16
Vx90 xm90 0 0
Gx90_1 x90 0 u1 0 1.15193289447181e-06
Rx91 x91 0 1
Fxc91_92 x91 0 Vx92 22093.311097251
Cx91 x91 xm91 1.91401504019507e-14
Vx91 xm91 0 0
Gx91_1 x91 0 u1 0 -4.26919507825896e-08
Rx92 x92 0 1
Fxc92_91 x92 0 Vx91 -39.79721599417
Cx92 x92 xm92 1.91401504019507e-14
Vx92 xm92 0 0
Gx92_1 x92 0 u1 0 1.6990207865072e-06
Rx93 x93 0 1
Fxc93_94 x93 0 Vx94 375.010594704786
Cx93 x93 xm93 2.78471100161717e-14
Vx93 xm93 0 0
Gx93_1 x93 0 u1 0 -6.39670943163263e-08
Rx94 x94 0 1
Fxc94_93 x94 0 Vx93 -1111.87956349289
Cx94 x94 xm94 2.78471100161717e-14
Vx94 xm94 0 0
Gx94_1 x94 0 u1 0 7.11237049063456e-05
Rx95 x95 0 1
Fxc95_96 x95 0 Vx96 13848.6792413956
Cx95 x95 xm95 7.87159377020613e-15
Vx95 xm95 0 0
Gx95_1 x95 0 u1 0 -3.19927800555257e-09
Rx96 x96 0 1
Fxc96_95 x96 0 Vx95 -371.264226747332
Cx96 x96 xm96 7.87159377020613e-15
Vx96 xm96 0 0
Gx96_1 x96 0 u1 0 1.18777747488122e-06
Rx97 x97 0 1
Fxc97_98 x97 0 Vx98 8.75011579927194
Cx97 x97 xm97 1.06813886291274e-12
Vx97 xm97 0 0
Gx97_1 x97 0 u1 0 -0.0406239272061045
Rx98 x98 0 1
Fxc98_97 x98 0 Vx97 -33.8662177042959
Cx98 x98 xm98 1.06813886291274e-12
Vx98 xm98 0 0
Gx98_1 x98 0 u1 0 1.37577876276541
Rx99 x99 0 1
Fxc99_100 x99 0 Vx100 10978.5499609988
Cx99 x99 xm99 5.25955260177112e-15
Vx99 xm99 0 0
Gx99_1 x99 0 u1 0 -1.85691748334487e-09
Rx100 x100 0 1
Fxc100_99 x100 0 Vx99 -1083.44784659305
Cx100 x100 xm100 5.25955260177112e-15
Vx100 xm100 0 0
Gx100_1 x100 0 u1 0 2.01187324863099e-06
Rx101 x101 0 1
Fxc101_102 x101 0 Vx102 628.943509862508
Cx101 x101 xm101 2.76085682247672e-14
Vx101 xm101 0 0
Gx101_1 x101 0 u1 0 -6.11681673256886e-08
Rx102 x102 0 1
Fxc102_101 x102 0 Vx101 -691.740691831882
Cx102 x102 xm102 2.76085682247672e-14
Vx102 xm102 0 0
Gx102_1 x102 0 u1 0 4.23125103839601e-05
Rx103 x103 0 1
Fxc103_104 x103 0 Vx104 606.599086946569
Cx103 x103 xm103 1.46519190092729e-14
Vx103 xm103 0 0
Gx103_1 x103 0 u1 0 -7.4927294404879e-09
Rx104 x104 0 1
Fxc104_103 x104 0 Vx103 -2562.99407233946
Cx104 x104 xm104 1.46519190092729e-14
Vx104 xm104 0 0
Gx104_1 x104 0 u1 0 1.92038211416139e-05
Rx105 x105 0 1
Fxc105_106 x105 0 Vx106 1463.83671763519
Cx105 x105 xm105 2.19788949285279e-14
Vx105 xm105 0 0
Gx105_1 x105 0 u1 0 -3.16477233836375e-08
Rx106 x106 0 1
Fxc106_105 x106 0 Vx105 -475.981534615473
Cx106 x106 xm106 2.19788949285279e-14
Vx106 xm106 0 0
Gx106_1 x106 0 u1 0 1.50637319432298e-05
Rx107 x107 0 1
Fxc107_108 x107 0 Vx108 511.712555444263
Cx107 x107 xm107 8.20375533487514e-14
Vx107 xm107 0 0
Gx107_1 x107 0 u1 0 -1.4465913024119e-06
Rx108 x108 0 1
Fxc108_107 x108 0 Vx107 -98.7065960828127
Cx108 x108 xm108 8.20375533487514e-14
Vx108 xm108 0 0
Gx108_1 x108 0 u1 0 0.000142788103384082
Rx109 x109 0 1
Fxc109_110 x109 0 Vx110 1840.08911733932
Cx109 x109 xm109 7.51272397073094e-15
Vx109 xm109 0 0
Gx109_1 x109 0 u1 0 -2.63856145339527e-09
Rx110 x110 0 1
Fxc110_109 x110 0 Vx109 -3281.78228604659
Cx110 x110 xm110 7.51272397073094e-15
Vx110 xm110 0 0
Gx110_1 x110 0 u1 0 8.65918423839794e-06
Rx111 x111 0 1
Fxc111_112 x111 0 Vx112 534.755990268543
Cx111 x111 xm111 1.25924088295157e-14
Vx111 xm111 0 0
Gx111_1 x111 0 u1 0 -2.0471663695567e-09
Rx112 x112 0 1
Fxc112_111 x112 0 Vx111 -4349.39000170155
Cx112 x112 xm112 1.25924088295157e-14
Vx112 xm112 0 0
Gx112_1 x112 0 u1 0 8.90392493956957e-06
Rx113 x113 0 1
Fxc113_114 x113 0 Vx114 149.866737948217
Cx113 x113 xm113 3.99671423619986e-14
Vx113 xm113 0 0
Gx113_1 x113 0 u1 0 -4.59375822675306e-08
Rx114 x114 0 1
Fxc114_113 x114 0 Vx113 -1531.92935076511
Cx114 x114 xm114 3.99671423619987e-14
Vx114 xm114 0 0
Gx114_1 x114 0 u1 0 7.03731305788168e-05
Rx115 x115 0 1
Fxc115_116 x115 0 Vx116 10545.6478758616
Cx115 x115 xm115 4.75295253243805e-15
Vx115 xm115 0 0
Gx115_1 x115 0 u1 0 -2.2487729127759e-09
Rx116 x116 0 1
Fxc116_115 x116 0 Vx115 -1448.25980659277
Cx116 x116 xm116 4.75295253243805e-15
Vx116 xm116 0 0
Gx116_1 x116 0 u1 0 3.25680742372789e-06
Rx117 x117 0 1
Fxc117_118 x117 0 Vx118 681.911447470694
Cx117 x117 xm117 3.41070990725561e-14
Vx117 xm117 0 0
Gx117_1 x117 0 u1 0 -7.94259015202656e-08
Rx118 x118 0 1
Fxc118_117 x118 0 Vx117 -437.145456629005
Cx118 x118 xm118 3.41070990725561e-14
Vx118 xm118 0 0
Gx118_1 x118 0 u1 0 3.47206719882468e-05
Rx119 x119 0 1
Fxc119_120 x119 0 Vx120 3927.86052023466
Cx119 x119 xm119 9.91623794270551e-15
Vx119 xm119 0 0
Gx119_1 x119 0 u1 0 -3.83159739907986e-09
Rx120 x120 0 1
Fxc120_119 x120 0 Vx119 -903.259681021793
Cx120 x120 xm120 9.91623794270551e-15
Vx120 xm120 0 0
Gx120_1 x120 0 u1 0 3.46092744449681e-06
Rx121 x121 0 1
Fxc121_122 x121 0 Vx122 672.490742606125
Cx121 x121 xm121 2.22232201775079e-14
Vx121 xm121 0 0
Gx121_1 x121 0 u1 0 -2.19041004489507e-08
Rx122 x122 0 1
Fxc122_121 x122 0 Vx121 -1093.78293184411
Cx122 x122 xm122 2.22232201775079e-14
Vx122 xm122 0 0
Gx122_1 x122 0 u1 0 2.39583312084613e-05
Rx123 x123 0 1
Fxc123_124 x123 0 Vx124 1424.64634121618
Cx123 x123 xm123 5.17797017606527e-15
Vx123 xm123 0 0
Gx123_1 x123 0 u1 0 -4.81135246026594e-10
Rx124 x124 0 1
Fxc124_123 x124 0 Vx123 -9202.05808625698
Cx124 x124 xm124 5.17797017606527e-15
Vx124 xm124 0 0
Gx124_1 x124 0 u1 0 4.42743448128226e-06
Rx125 x125 0 1
Fxc125_126 x125 0 Vx126 393.964226248637
Cx125 x125 xm125 4.46596707298567e-14
Vx125 xm125 0 0
Gx125_1 x125 0 u1 0 -2.47449617543097e-07
Rx126 x126 0 1
Fxc126_125 x126 0 Vx125 -453.75387202112
Cx126 x126 xm126 4.46596707298567e-14
Vx126 xm126 0 0
Gx126_1 x126 0 u1 0 0.000112281222090325
Rx127 x127 0 1
Fxc127_128 x127 0 Vx128 1174.69871746606
Cx127 x127 xm127 1.25147099405371e-14
Vx127 xm127 0 0
Gx127_1 x127 0 u1 0 -6.77009308214809e-09
Rx128 x128 0 1
Fxc128_127 x128 0 Vx127 -1964.69277457512
Cx128 x128 xm128 1.25147099405371e-14
Vx128 xm128 0 0
Gx128_1 x128 0 u1 0 1.33011529616974e-05
Rx129 x129 0 1
Fxc129_130 x129 0 Vx130 1415.58288437931
Cx129 x129 xm129 3.07868023406084e-14
Vx129 xm129 0 0
Gx129_1 x129 0 u1 0 -1.0579300204017e-07
Rx130 x130 0 1
Fxc130_129 x130 0 Vx129 -267.277316448364
Cx130 x130 xm130 3.07868023406084e-14
Vx130 xm130 0 0
Gx130_1 x130 0 u1 0 2.8276069684313e-05
Rx131 x131 0 1
Fxc131_132 x131 0 Vx132 805.91935992515
Cx131 x131 xm131 5.4585280782342e-15
Vx131 xm131 0 0
Gx131_1 x131 0 u1 0 -5.60153059722672e-10
Rx132 x132 0 1
Fxc132_131 x132 0 Vx131 -14854.0843048736
Cx132 x132 xm132 5.4585280782342e-15
Vx132 xm132 0 0
Gx132_1 x132 0 u1 0 8.32056077275346e-06
Rx133 x133 0 1
Fxc133_134 x133 0 Vx134 12.6887732169287
Cx133 x133 xm133 2.51329289587019e-12
Vx133 xm133 0 0
Gx133_1 x133 0 u1 0 -1.07071429988905
Rx134 x134 0 1
Fxc134_133 x134 0 Vx133 -5.34166240603459
Cx134 x134 xm134 2.51329289587019e-12
Vx134 xm134 0 0
Gx134_1 x134 0 u1 0 5.71939432332099
Rx135 x135 0 1
Fxc135_136 x135 0 Vx136 135.73862234201
Cx135 x135 xm135 3.57049647256315e-13
Vx135 xm135 0 0
Gx135_1 x135 0 u1 0 -0.000179883802904531
Rx136 x136 0 1
Fxc136_135 x136 0 Vx135 -23.7418745932653
Cx136 x136 xm136 3.57049647256315e-13
Vx136 xm136 0 0
Gx136_1 x136 0 u1 0 0.00427077868991902
Rx137 x137 0 1
Fxc137_138 x137 0 Vx138 428.13489270737
Cx137 x137 xm137 4.5035441503013e-14
Vx137 xm137 0 0
Gx137_1 x137 0 u1 0 -1.37186306748478e-07
Rx138 x138 0 1
Fxc138_137 x138 0 Vx137 -427.576045386489
Cx138 x138 xm138 4.5035441503013e-14
Vx138 xm138 0 0
Gx138_1 x138 0 u1 0 5.86575785206919e-05
Rx139 x139 0 1
Fxc139_140 x139 0 Vx140 1535.85616609788
Cx139 x139 xm139 8.56467633357547e-15
Vx139 xm139 0 0
Gx139_1 x139 0 u1 0 -1.22149616518128e-09
Rx140 x140 0 1
Fxc140_139 x140 0 Vx139 -3327.27372575882
Cx140 x140 xm140 8.56467633357547e-15
Vx140 xm140 0 0
Gx140_1 x140 0 u1 0 4.06425209652283e-06
Rx141 x141 0 1
Fxc141_142 x141 0 Vx142 171.094267029573
Cx141 x141 xm141 8.27372304605411e-14
Vx141 xm141 0 0
Gx141_1 x141 0 u1 0 -5.0313737612082e-07
Rx142 x142 0 1
Fxc142_141 x142 0 Vx141 -343.938297227506
Cx142 x142 xm142 8.27372304605411e-14
Vx142 xm142 0 0
Gx142_1 x142 0 u1 0 0.00017304821241451
Rx143 x143 0 1
Fxc143_144 x143 0 Vx144 1206.58470663483
Cx143 x143 xm143 1.66721817308413e-14
Vx143 xm143 0 0
Gx143_1 x143 0 u1 0 -1.35794105530886e-08
Rx144 x144 0 1
Fxc144_143 x144 0 Vx143 -1123.56307144083
Cx144 x144 xm144 1.66721817308413e-14
Vx144 xm144 0 0
Gx144_1 x144 0 u1 0 1.52573242293843e-05
Rx145 x145 0 1
Fxc145_146 x145 0 Vx146 2195.49276741284
Cx145 x145 xm145 7.00529634671639e-14
Vx145 xm145 0 0
Gx145_1 x145 0 u1 0 -9.28851351565625e-07
Rx146 x146 0 1
Fxc146_145 x146 0 Vx145 -35.0443706113712
Cx146 x146 xm146 7.0052963467164e-14
Vx146 xm146 0 0
Gx146_1 x146 0 u1 0 3.25510110071388e-05
Rx147 x147 0 1
Fxc147_148 x147 0 Vx148 17296.6665638803
Cx147 x147 xm147 1.10677227211622e-16
Vx147 xm147 0 0
Gx147_1 x147 0 u1 0 -8.89803244945423e-13
Rx148 x148 0 1
Fxc148_147 x148 0 Vx147 -1895934.61538509
Cx148 x148 xm148 1.10677227211622e-16
Vx148 xm148 0 0
Gx148_1 x148 0 u1 0 1.687008772974e-06
Rx149 x149 0 1
Fxc149_150 x149 0 Vx150 9028.42462041655
Cx149 x149 xm149 1.5846769699005e-14
Vx149 xm149 0 0
Gx149_1 x149 0 u1 0 -1.03467434743729e-08
Rx150 x150 0 1
Fxc150_149 x150 0 Vx149 -175.300173553119
Cx150 x150 xm150 1.5846769699005e-14
Vx150 xm150 0 0
Gx150_1 x150 0 u1 0 1.81378592676718e-06
Rx151 x151 0 1
Fxc151_152 x151 0 Vx152 755.243881753823
Cx151 x151 xm151 4.12031373830175e-14
Vx151 xm151 0 0
Gx151_1 x151 0 u1 0 -3.36445271183827e-07
Rx152 x152 0 1
Fxc152_151 x152 0 Vx151 -300.360256673079
Cx152 x152 xm152 4.12031373830175e-14
Vx152 xm152 0 0
Gx152_1 x152 0 u1 0 0.000101054788009218
Rx153 x153 0 1
Fxc153_154 x153 0 Vx154 2072.1952183899
Cx153 x153 xm153 1.43266280058829e-14
Vx153 xm153 0 0
Gx153_1 x153 0 u1 0 -9.98194844813138e-09
Rx154 x154 0 1
Fxc154_153 x154 0 Vx153 -900.3118843563
Cx154 x154 xm154 1.43266280058829e-14
Vx154 xm154 0 0
Gx154_1 x154 0 u1 0 8.98686681688461e-06
Rx155 x155 0 1
Fxc155_156 x155 0 Vx156 358.087520404934
Cx155 x155 xm155 9.37589835741656e-14
Vx155 xm155 0 0
Gx155_1 x155 0 u1 0 -2.92937751883025e-06
Rx156 x156 0 1
Fxc156_155 x156 0 Vx155 -123.239388501282
Cx156 x156 xm156 9.37589835741656e-14
Vx156 xm156 0 0
Gx156_1 x156 0 u1 0 0.000361014694110043
Rx157 x157 0 1
Fxc157_158 x157 0 Vx158 548.100843242006
Cx157 x157 xm157 2.94431934184726e-15
Vx157 xm157 0 0
Gx157_1 x157 0 u1 0 -4.42823423287936e-11
Rx158 x158 0 1
Fxc158_157 x158 0 Vx157 -82185.5234858855
Cx158 x158 xm158 2.94431934184726e-15
Vx158 xm158 0 0
Gx158_1 x158 0 u1 0 3.63936748547309e-06
Rx159 x159 0 1
Fxc159_160 x159 0 Vx160 790212.37398732
Cx159 x159 xm159 1.38008738267159e-16
Vx159 xm159 0 0
Gx159_1 x159 0 u1 0 -2.79862793496414e-12
Rx160 x160 0 1
Fxc160_159 x160 0 Vx159 -26176.8898998116
Cx160 x160 xm160 1.38008738267159e-16
Vx160 xm160 0 0
Gx160_1 x160 0 u1 0 7.32593753240934e-08
Rx161 x161 0 1
Fxc161_162 x161 0 Vx162 143.767839089496
Cx161 x161 xm161 3.31616743972311e-14
Vx161 xm161 0 0
Gx161_1 x161 0 u1 0 -4.95582337534821e-08
Rx162 x162 0 1
Fxc162_161 x162 0 Vx161 -2445.85926995736
Cx162 x162 xm162 3.31616743972311e-14
Vx162 xm162 0 0
Gx162_1 x162 0 u1 0 0.000121212465428668
Rx163 x163 0 1
Fxc163_164 x163 0 Vx164 32.1947548695074
Cx163 x163 xm163 6.8171023360865e-13
Vx163 xm163 0 0
Gx163_1 x163 0 u1 0 -0.00425318185303686
Rx164 x164 0 1
Fxc164_163 x164 0 Vx163 -28.9379488109184
Cx164 x164 xm164 6.8171023360865e-13
Vx164 xm164 0 0
Gx164_1 x164 0 u1 0 0.123078358746708
Rx165 x165 0 1
Fxc165_166 x165 0 Vx166 10560.8526810331
Cx165 x165 xm165 1.6412792293327e-15
Vx165 xm165 0 0
Gx165_1 x165 0 u1 0 -2.32902315011842e-10
Rx166 x166 0 1
Fxc166_165 x166 0 Vx165 -14286.9129172589
Cx166 x166 xm166 1.6412792293327e-15
Vx166 xm166 0 0
Gx166_1 x166 0 u1 0 3.32745509280219e-06
Rx167 x167 0 1
Fxc167_168 x167 0 Vx168 68.448808395086
Cx167 x167 xm167 2.0277279276718e-14
Vx167 xm167 0 0
Gx167_1 x167 0 u1 0 -1.21053960220682e-09
Rx168 x168 0 1
Fxc168_167 x168 0 Vx167 -15513.1812004414
Cx168 x168 xm168 2.0277279276718e-14
Vx168 xm168 0 0
Gx168_1 x168 0 u1 0 1.87793201993446e-05
Rx169 x169 0 1
Fxc169_170 x169 0 Vx170 1487.45510739481
Cx169 x169 xm169 9.54778893264496e-15
Vx169 xm169 0 0
Gx169_1 x169 0 u1 0 -1.50371032679042e-09
Rx170 x170 0 1
Fxc170_169 x170 0 Vx169 -3012.21772107701
Cx170 x170 xm170 9.54778893264496e-15
Vx170 xm170 0 0
Gx170_1 x170 0 u1 0 4.5295028937246e-06
Rx171 x171 0 1
Fxc171_172 x171 0 Vx172 2121.83105981255
Cx171 x171 xm171 1.33797401275805e-14
Vx171 xm171 0 0
Gx171_1 x171 0 u1 0 -4.60700732431939e-09
Rx172 x172 0 1
Fxc172_171 x172 0 Vx171 -1085.31420689364
Cx172 x172 xm172 1.33797401275805e-14
Vx172 xm172 0 0
Gx172_1 x172 0 u1 0 5.00005050034689e-06
Rx173 x173 0 1
Fxc173_174 x173 0 Vx174 67595.9477186301
Cx173 x173 xm173 8.17600979330828e-15
Vx173 xm173 0 0
Gx173_1 x173 0 u1 0 -1.74203636305824e-09
Rx174 x174 0 1
Fxc174_173 x174 0 Vx173 -92.636632352269
Cx174 x174 xm174 8.17600979330828e-15
Vx174 xm174 0 0
Gx174_1 x174 0 u1 0 1.6137638210891e-07
Rx175 x175 0 1
Fxc175_176 x175 0 Vx176 1294.86265829018
Cx175 x175 xm175 1.96425850879399e-14
Vx175 xm175 0 0
Gx175_1 x175 0 u1 0 -1.12401587857913e-08
Rx176 x176 0 1
Fxc176_175 x176 0 Vx175 -862.960806550733
Cx176 x176 xm176 1.96425850879399e-14
Vx176 xm176 0 0
Gx176_1 x176 0 u1 0 9.69981649154475e-06
Rx177 x177 0 1
Fxc177_178 x177 0 Vx178 665.831950219072
Cx177 x177 xm177 1.88286053329382e-14
Vx177 xm177 0 0
Gx177_1 x177 0 u1 0 -8.58590225617211e-09
Rx178 x178 0 1
Fxc178_177 x178 0 Vx177 -1842.34892403804
Cx178 x178 xm178 1.88286053329382e-14
Vx178 xm178 0 0
Gx178_1 x178 0 u1 0 1.58182277835544e-05
Rx179 x179 0 1
Fxc179_180 x179 0 Vx180 2107.82872048532
Cx179 x179 xm179 1.88018559993273e-14
Vx179 xm179 0 0
Gx179_1 x179 0 u1 0 -1.3085235693506e-08
Rx180 x180 0 1
Fxc180_179 x180 0 Vx179 -573.89097712545
Cx180 x180 xm180 1.88018559993273e-14
Vx180 xm180 0 0
Gx180_1 x180 0 u1 0 7.509498698063e-06
Rx181 x181 0 1
Fxc181_182 x181 0 Vx182 145368.494187308
Cx181 x181 xm181 1.24637336182943e-15
Vx181 xm181 0 0
Gx181_1 x181 0 u1 0 -1.53914135759411e-10
Rx182 x182 0 1
Fxc182_181 x182 0 Vx181 -1844.10849027669
Cx182 x182 xm182 1.24637336182943e-15
Vx182 xm182 0 0
Gx182_1 x182 0 u1 0 2.83834364527529e-07
Rx183 x183 0 1
Fxc183_184 x183 0 Vx184 1093.45177134477
Cx183 x183 xm183 9.701039005748e-15
Vx183 xm183 0 0
Gx183_1 x183 0 u1 0 -1.65742015547723e-09
Rx184 x184 0 1
Fxc184_183 x184 0 Vx183 -4102.13224941861
Cx184 x184 xm184 9.701039005748e-15
Vx184 xm184 0 0
Gx184_1 x184 0 u1 0 6.79895667061955e-06
Rx185 x185 0 1
Fxc185_186 x185 0 Vx186 523.771889282841
Cx185 x185 xm185 2.77515669599418e-14
Vx185 xm185 0 0
Gx185_1 x185 0 u1 0 -2.22678753339474e-08
Rx186 x186 0 1
Fxc186_185 x186 0 Vx185 -1052.54221731094
Cx186 x186 xm186 2.77515669599418e-14
Vx186 xm186 0 0
Gx186_1 x186 0 u1 0 2.34378788787966e-05
Rx187 x187 0 1
Fxc187_188 x187 0 Vx188 58.1057285274661
Cx187 x187 xm187 1.90385021922328e-12
Vx187 xm187 0 0
Gx187_1 x187 0 u1 0 -0.334532302795897
Rx188 x188 0 1
Fxc188_187 x188 0 Vx187 -2.25235219973742
Cx188 x188 xm188 1.90385021922328e-12
Vx188 xm188 0 0
Gx188_1 x188 0 u1 0 0.753484568085563
Rx189 x189 0 1
Fxc189_190 x189 0 Vx190 219.689439110443
Cx189 x189 xm189 4.13080608699608e-13
Vx189 xm189 0 0
Gx189_1 x189 0 u1 0 -0.000913721674204237
Rx190 x190 0 1
Fxc190_189 x190 0 Vx189 -12.557817545699
Cx190 x190 xm190 4.13080608699608e-13
Vx190 xm190 0 0
Gx190_1 x190 0 u1 0 0.0114743500722075
Rx191 x191 0 1
Fxc191_192 x191 0 Vx192 17.1225668717222
Cx191 x191 xm191 3.88335929258945e-13
Vx191 xm191 0 0
Gx191_1 x191 0 u1 0 -0.000489166922433175
Rx192 x192 0 1
Fxc192_191 x192 0 Vx191 -177.554997252642
Cx192 x192 xm192 3.88335929258945e-13
Vx192 xm192 0 0
Gx192_1 x192 0 u1 0 0.0868540315687058
Rx193 x193 0 1
Fxc193_194 x193 0 Vx194 130.665838089954
Cx193 x193 xm193 2.37282917151686e-13
Vx193 xm193 0 0
Gx193_1 x193 0 u1 0 -0.000129064393457941
Rx194 x194 0 1
Fxc194_193 x194 0 Vx193 -61.8972239115515
Cx194 x194 xm194 2.37282917151686e-13
Vx194 xm194 0 0
Gx194_1 x194 0 u1 0 0.00798872766087474
Rx195 x195 0 1
Fxc195_196 x195 0 Vx196 312.778730468328
Cx195 x195 xm195 1.91607970073068e-14
Vx195 xm195 0 0
Gx195_1 x195 0 u1 0 -3.36657106871807e-09
Rx196 x196 0 1
Fxc196_195 x196 0 Vx195 -3862.43333752286
Cx196 x196 xm196 1.91607970073068e-14
Vx196 xm196 0 0
Gx196_1 x196 0 u1 0 1.30031563289567e-05
Rx197 x197 0 1
Fxc197_198 x197 0 Vx198 5980.89782530992
Cx197 x197 xm197 2.33334731840831e-14
Vx197 xm197 0 0
Gx197_1 x197 0 u1 0 -2.61960376680653e-08
Rx198 x198 0 1
Fxc198_197 x198 0 Vx197 -143.386988081432
Cx198 x198 xm198 2.33334731840831e-14
Vx198 xm198 0 0
Gx198_1 x198 0 u1 0 3.75617094089162e-06
Rx199 x199 0 1
Fxc199_200 x199 0 Vx200 17303.952214653
Cx199 x199 xm199 2.2448315996525e-14
Vx199 xm199 0 0
Gx199_1 x199 0 u1 0 -2.61530019384294e-08
Rx200 x200 0 1
Fxc200_199 x200 0 Vx199 -53.2750828597523
Cx200 x200 xm200 2.2448315996525e-14
Vx200 xm200 0 0
Gx200_1 x200 0 u1 0 1.39330334530109e-06
Rx201 x201 0 1
Fxc201_202 x201 0 Vx202 651.819322179663
Cx201 x201 xm201 5.50128571655933e-15
Vx201 xm201 0 0
Gx201_1 x201 0 u1 0 -1.2592688608217e-10
Rx202 x202 0 1
Fxc202_201 x202 0 Vx201 -23353.9097719269
Cx202 x202 xm202 5.50128571655933e-15
Vx202 xm202 0 0
Gx202_1 x202 0 u1 0 2.9408851354227e-06
Rx203 x203 0 1
Fxc203_204 x203 0 Vx204 442.050502332637
Cx203 x203 xm203 5.82585824065102e-14
Vx203 xm203 0 0
Gx203_1 x203 0 u1 0 -2.92422788971848e-07
Rx204 x204 0 1
Fxc204_203 x204 0 Vx203 -301.790448356168
Cx204 x204 xm204 5.82585824065102e-14
Vx204 xm204 0 0
Gx204_1 x204 0 u1 0 8.82504045933753e-05
Rx205 x205 0 1
Fxc205_206 x205 0 Vx206 2998.89025351833
Cx205 x205 xm205 4.64126067377759e-16
Vx205 xm205 0 0
Gx205_1 x205 0 u1 0 -2.86192572243224e-12
Rx206 x206 0 1
Fxc206_205 x206 0 Vx205 -699177.783986947
Cx206 x206 xm206 4.64126067377759e-16
Vx206 xm206 0 0
Gx206_1 x206 0 u1 0 2.00099488454542e-06
Rx207 x207 0 1
Fxc207_208 x207 0 Vx208 67732.5032338237
Cx207 x207 xm207 4.79316217773287e-15
Vx207 xm207 0 0
Gx207_1 x207 0 u1 0 -6.73420852715933e-10
Rx208 x208 0 1
Fxc208_207 x208 0 Vx207 -287.163158878416
Cx208 x208 xm208 4.79316217773287e-15
Vx208 xm208 0 0
Gx208_1 x208 0 u1 0 1.93381659320504e-07
Rx209 x209 0 1
Fxc209_210 x209 0 Vx210 3.01827543424663
Cx209 x209 xm209 4.88202959865766e-12
Vx209 xm209 0 0
Gx209_1 x209 0 u1 0 -0.580994809682523
Rx210 x210 0 1
Fxc210_209 x210 0 Vx209 -8.07020945616114
Cx210 x210 xm210 4.88202959865766e-12
Vx210 xm210 0 0
Gx210_1 x210 0 u1 0 4.68874980708043
Rx211 x211 0 1
Fxc211_212 x211 0 Vx212 4564.13733356228
Cx211 x211 xm211 3.10944035248846e-15
Vx211 xm211 0 0
Gx211_1 x211 0 u1 0 -3.80020778736851e-11
Rx212 x212 0 1
Fxc212_211 x212 0 Vx211 -10739.8654828533
Cx212 x212 xm212 3.10944035248846e-15
Vx212 xm212 0 0
Gx212_1 x212 0 u1 0 4.08137204432294e-07
Rx213 x213 0 1
Fxc213_214 x213 0 Vx214 1037.6188837696
Cx213 x213 xm213 2.0409012950473e-14
Vx213 xm213 0 0
Gx213_1 x213 0 u1 0 -1.55099419235932e-08
Rx214 x214 0 1
Fxc214_213 x214 0 Vx213 -1108.00286318647
Cx214 x214 xm214 2.0409012950473e-14
Vx214 xm214 0 0
Gx214_1 x214 0 u1 0 1.71850600591971e-05
Rx215 x215 0 1
Fxc215_216 x215 0 Vx216 804.603657950695
Cx215 x215 xm215 4.35243189785395e-14
Vx215 xm215 0 0
Gx215_1 x215 0 u1 0 -3.06722495558031e-07
Rx216 x216 0 1
Fxc216_215 x216 0 Vx215 -317.118282736887
Cx216 x216 xm216 4.35243189785395e-14
Vx216 xm216 0 0
Gx216_1 x216 0 u1 0 9.72673110681353e-05
Rx217 x217 0 1
Fxc217_218 x217 0 Vx218 608.839969558945
Cx217 x217 xm217 4.3066796599514e-14
Vx217 xm217 0 0
Gx217_1 x217 0 u1 0 -2.4503725635058e-07
Rx218 x218 0 1
Fxc218_217 x218 0 Vx217 -426.4477553338
Cx218 x218 xm218 4.30667965995139e-14
Vx218 xm218 0 0
Gx218_1 x218 0 u1 0 0.000104495587943858
Rx219 x219 0 1
Fxc219_220 x219 0 Vx220 452.38998904912
Cx219 x219 xm219 3.11541373257599e-14
Vx219 xm219 0 0
Gx219_1 x219 0 u1 0 -4.08592970341204e-08
Rx220 x220 0 1
Fxc220_219 x220 0 Vx219 -1106.24273199186
Cx220 x220 xm220 3.11541373257599e-14
Vx220 xm220 0 0
Gx220_1 x220 0 u1 0 4.52003003782921e-05
Rx221 x221 0 1
Fxc221_222 x221 0 Vx222 55.0743971075051
Cx221 x221 xm221 1.22063164496342e-13
Vx221 xm221 0 0
Gx221_1 x221 0 u1 0 -9.05490804118085e-07
Rx222 x222 0 1
Fxc222_221 x222 0 Vx221 -606.919557716483
Cx222 x222 xm222 1.22063164496342e-13
Vx222 xm222 0 0
Gx222_1 x222 0 u1 0 0.000549560078351691
Rx223 x223 0 1
Fxc223_224 x223 0 Vx224 45.0132851649246
Cx223 x223 xm223 2.56056905033321e-14
Vx223 xm223 0 0
Gx223_1 x223 0 u1 0 -1.78203953081713e-09
Rx224 x224 0 1
Fxc224_223 x224 0 Vx223 -16641.7038077781
Cx224 x224 xm224 2.56056905033321e-14
Vx224 xm224 0 0
Gx224_1 x224 0 u1 0 2.96561740456104e-05
Rx225 x225 0 1
Fxc225_226 x225 0 Vx226 634.572639152941
Cx225 x225 xm225 9.10350048138882e-15
Vx225 xm225 0 0
Gx225_1 x225 0 u1 0 -1.95448277992277e-10
Rx226 x226 0 1
Fxc226_225 x226 0 Vx225 -9800.48029981583
Cx226 x226 xm226 9.10350048138882e-15
Vx226 xm226 0 0
Gx226_1 x226 0 u1 0 1.91548699809624e-06
Rx227 x227 0 1
Fxc227_228 x227 0 Vx228 1040.01664265881
Cx227 x227 xm227 1.25795884003576e-14
Vx227 xm227 0 0
Gx227_1 x227 0 u1 0 -3.67639423457434e-09
Rx228 x228 0 1
Fxc228_227 x228 0 Vx227 -3002.37874781419
Cx228 x228 xm228 1.25795884003576e-14
Vx228 xm228 0 0
Gx228_1 x228 0 u1 0 1.10379279184726e-05
Rx229 x229 0 1
Fxc229_230 x229 0 Vx230 16331.7452099969
Cx229 x229 xm229 6.42832682389733e-15
Vx229 xm229 0 0
Gx229_1 x229 0 u1 0 -7.56666790105865e-10
Rx230 x230 0 1
Fxc230_229 x230 0 Vx229 -751.765722658087
Cx230 x230 xm230 6.42832682389733e-15
Vx230 xm230 0 0
Gx230_1 x230 0 u1 0 5.68836156275311e-07
Rx231 x231 0 1
Fxc231_232 x231 0 Vx232 269.115226072413
Cx231 x231 xm231 3.78461462762688e-14
Vx231 xm231 0 0
Gx231_1 x231 0 u1 0 -1.76404608106008e-08
Rx232 x232 0 1
Fxc232_231 x232 0 Vx231 -1333.12202322767
Cx232 x232 xm232 3.78461462762688e-14
Vx232 xm232 0 0
Gx232_1 x232 0 u1 0 2.35168868064965e-05
Rx233 x233 0 1
Fxc233_234 x233 0 Vx234 10614.3274520747
Cx233 x233 xm233 7.47163154472277e-15
Vx233 xm233 0 0
Gx233_1 x233 0 u1 0 -3.61593102718078e-09
Rx234 x234 0 1
Fxc234_233 x234 0 Vx233 -846.415172955531
Cx234 x234 xm234 7.47163154472277e-15
Vx234 xm234 0 0
Gx234_1 x234 0 u1 0 3.06057888576649e-06
Rx235 x235 0 1
Fxc235_236 x235 0 Vx236 9390.43673298885
Cx235 x235 xm235 4.17550450563194e-14
Vx235 xm235 0 0
Gx235_1 x235 0 u1 0 -1.47268138397953e-07
Rx236 x236 0 1
Fxc236_235 x236 0 Vx235 -30.6038047151082
Cx236 x236 xm236 4.17550450563194e-14
Vx236 xm236 0 0
Gx236_1 x236 0 u1 0 4.50696534828848e-06
Rx237 x237 0 1
Fxc237_238 x237 0 Vx238 545.751476568648
Cx237 x237 xm237 3.5696335326637e-13
Vx237 xm237 0 0
Gx237_1 x237 0 u1 0 -6.27738180736851e-05
Rx238 x238 0 1
Fxc238_237 x238 0 Vx237 -7.72133018190495
Cx238 x238 xm238 3.5696335326637e-13
Vx238 xm238 0 0
Gx238_1 x238 0 u1 0 0.000484697376125755
Rx239 x239 0 1
Fxc239_240 x239 0 Vx240 830.303215997316
Cx239 x239 xm239 1.92605907935797e-14
Vx239 xm239 0 0
Gx239_1 x239 0 u1 0 -7.31844571930659e-09
Rx240 x240 0 1
Fxc240_239 x240 0 Vx239 -1692.85982852407
Cx240 x240 xm240 1.92605907935797e-14
Vx240 xm240 0 0
Gx240_1 x240 0 u1 0 1.23891027654481e-05
Rx241 x241 0 1
Fxc241_242 x241 0 Vx242 1744.54142376656
Cx241 x241 xm241 4.96085474377487e-14
Vx241 xm241 0 0
Gx241_1 x241 0 u1 0 -1.35906058097832e-07
Rx242 x242 0 1
Fxc242_241 x242 0 Vx241 -121.977780367775
Cx242 x242 xm242 4.96085474377487e-14
Vx242 xm242 0 0
Gx242_1 x242 0 u1 0 1.65775193053074e-05
Rx243 x243 0 1
Fxc243_244 x243 0 Vx244 3634.98988839577
Cx243 x243 xm243 1.34382674878936e-14
Vx243 xm243 0 0
Gx243_1 x243 0 u1 0 -5.54834431265805e-09
Rx244 x244 0 1
Fxc244_243 x244 0 Vx243 -802.443381508567
Cx244 x244 xm244 1.34382674878936e-14
Vx244 xm244 0 0
Gx244_1 x244 0 u1 0 4.45223217202315e-06
Rx245 x245 0 1
Fxc245_246 x245 0 Vx246 449.441625819739
Cx245 x245 xm245 8.72908617003218e-15
Vx245 xm245 0 0
Gx245_1 x245 0 u1 0 -1.27030558275292e-10
Rx246 x246 0 1
Fxc246_245 x246 0 Vx245 -15597.8330576724
Cx246 x246 xm246 8.72908617003218e-15
Vx246 xm246 0 0
Gx246_1 x246 0 u1 0 1.98140144120094e-06
Rx247 x247 0 1
Fxc247_248 x247 0 Vx248 828.634673955662
Cx247 x247 xm247 1.41656257366965e-14
Vx247 xm247 0 0
Gx247_1 x247 0 u1 0 -2.36298078557977e-09
Rx248 x248 0 1
Fxc248_247 x248 0 Vx247 -3234.52262828574
Cx248 x248 xm248 1.41656257366965e-14
Vx248 xm248 0 0
Gx248_1 x248 0 u1 0 7.64311482116218e-06
Rx249 x249 0 1
Fxc249_250 x249 0 Vx250 32.8102482604173
Cx249 x249 xm249 6.46803689263805e-13
Vx249 xm249 0 0
Gx249_1 x249 0 u1 0 -0.000306808352885927
Rx250 x250 0 1
Fxc250_249 x250 0 Vx249 -42.2128957593941
Cx250 x250 xm250 6.46803689263805e-13
Vx250 xm250 0 0
Gx250_1 x250 0 u1 0 0.012951269018485
Rx251 x251 0 1
Fxc251_252 x251 0 Vx252 20.7159804395296
Cx251 x251 xm251 2.59067693849385e-14
Vx251 xm251 0 0
Gx251_1 x251 0 u1 0 -5.4103932488581e-10
Rx252 x252 0 1
Fxc252_251 x252 0 Vx251 -39006.7874393571
Cx252 x252 xm252 2.59067693849385e-14
Vx252 xm252 0 0
Gx252_1 x252 0 u1 0 2.11042059421541e-05
Rx253 x253 0 1
Fxc253_254 x253 0 Vx254 55476.2121981388
Cx253 x253 xm253 3.81925234457657e-15
Vx253 xm253 0 0
Gx253_1 x253 0 u1 0 -1.33679062639461e-09
Rx254 x254 0 1
Fxc254_253 x254 0 Vx253 -676.974225594198
Cx254 x254 xm254 3.81925234457657e-15
Vx254 xm254 0 0
Gx254_1 x254 0 u1 0 9.04972799085073e-07
Rx255 x255 0 1
Fxc255_256 x255 0 Vx256 97.0295254717883
Cx255 x255 xm255 5.61704850831073e-14
Vx255 xm255 0 0
Gx255_1 x255 0 u1 0 -5.8424974974284e-08
Rx256 x256 0 1
Fxc256_255 x256 0 Vx255 -1811.31547032578
Cx256 x256 xm256 5.61704850831073e-14
Vx256 xm256 0 0
Gx256_1 x256 0 u1 0 0.000105826061024317
Rx257 x257 0 1
Fxc257_258 x257 0 Vx258 502.936111839346
Cx257 x257 xm257 4.39028211648867e-14
Vx257 xm257 0 0
Gx257_1 x257 0 u1 0 -1.04815843750513e-07
Rx258 x258 0 1
Fxc258_257 x258 0 Vx257 -574.814159191333
Cx258 x258 xm258 4.39028211648867e-14
Vx258 xm258 0 0
Gx258_1 x258 0 u1 0 6.02496310953811e-05
Rx259 x259 0 1
Fxc259_260 x259 0 Vx260 340.212991165746
Cx259 x259 xm259 3.387890067806e-14
Vx259 xm259 0 0
Gx259_1 x259 0 u1 0 -2.99261508839012e-08
Rx260 x260 0 1
Fxc260_259 x260 0 Vx259 -1438.82674069849
Cx260 x260 xm260 3.387890067806e-14
Vx260 xm260 0 0
Gx260_1 x260 0 u1 0 4.30585461379349e-05
Rx261 x261 0 1
Fxc261_262 x261 0 Vx262 6140.96620508896
Cx261 x261 xm261 2.71987544670807e-14
Vx261 xm261 0 0
Gx261_1 x261 0 u1 0 -5.15494367597002e-08
Rx262 x262 0 1
Fxc262_261 x262 0 Vx261 -124.526326417509
Cx262 x262 xm262 2.71987544670807e-14
Vx262 xm262 0 0
Gx262_1 x262 0 u1 0 6.41926198857718e-06
Rx263 x263 0 1
Fxc263_264 x263 0 Vx264 23.2258235715275
Cx263 x263 xm263 9.59156105724643e-14
Vx263 xm263 0 0
Gx263_1 x263 0 u1 0 -1.93889616268584e-07
Rx264 x264 0 1
Fxc264_263 x264 0 Vx263 -2661.08512464258
Cx264 x264 xm264 9.59156105724643e-14
Vx264 xm264 0 0
Gx264_1 x264 0 u1 0 0.000515956773674987
Rx265 x265 0 1
Fxc265_266 x265 0 Vx266 6037.59308361684
Cx265 x265 xm265 2.29533381547327e-14
Vx265 xm265 0 0
Gx265_1 x265 0 u1 0 -7.20917175970576e-08
Rx266 x266 0 1
Fxc266_265 x266 0 Vx265 -179.685592173743
Cx266 x266 xm266 2.29533381547327e-14
Vx266 xm266 0 0
Gx266_1 x266 0 u1 0 1.29538429672496e-05
Rx267 x267 0 1
Fxc267_268 x267 0 Vx268 1723.34134129715
Cx267 x267 xm267 4.98360784941284e-15
Vx267 xm267 0 0
Gx267_1 x267 0 u1 0 -1.28100890992794e-09
Rx268 x268 0 1
Fxc268_267 x268 0 Vx267 -13376.4383111057
Cx268 x268 xm268 4.98360784941284e-15
Vx268 xm268 0 0
Gx268_1 x268 0 u1 0 1.71353366596279e-05
Rx269 x269 0 1
Fxc269_270 x269 0 Vx270 1946.83794295379
Cx269 x269 xm269 2.42570294480808e-15
Vx269 xm269 0 0
Gx269_1 x269 0 u1 0 -1.14736422852399e-10
Rx270 x270 0 1
Fxc270_269 x270 0 Vx269 -50738.1413317836
Cx270 x270 xm270 2.42570294480808e-15
Vx270 xm270 0 0
Gx270_1 x270 0 u1 0 5.82151283858828e-06
Rx271 x271 0 1
Fxc271_272 x271 0 Vx272 134853.780166479
Cx271 x271 xm271 2.25473411609031e-15
Vx271 xm271 0 0
Gx271_1 x271 0 u1 0 -2.23100402651917e-10
Rx272 x272 0 1
Fxc272_271 x272 0 Vx271 -853.695796444358
Cx272 x272 xm272 2.25473411609031e-15
Vx272 xm272 0 0
Gx272_1 x272 0 u1 0 1.90459875928985e-07
Rx273 x273 0 1
Fxc273_274 x273 0 Vx274 1089.95157450767
Cx273 x273 xm273 1.48732812338964e-14
Vx273 xm273 0 0
Gx273_1 x273 0 u1 0 -2.43574581796807e-09
Rx274 x274 0 1
Fxc274_273 x274 0 Vx273 -2445.71612398201
Cx274 x274 xm274 1.48732812338964e-14
Vx274 xm274 0 0
Gx274_1 x274 0 u1 0 5.95714282092626e-06
Rx275 x275 0 1
Fxc275_276 x275 0 Vx276 4228.87990000677
Cx275 x275 xm275 5.99616853581674e-15
Vx275 xm275 0 0
Gx275_1 x275 0 u1 0 -6.48417207466053e-10
Rx276 x276 0 1
Fxc276_275 x276 0 Vx275 -3927.08321264857
Cx276 x276 xm276 5.99616853581674e-15
Vx276 xm276 0 0
Gx276_1 x276 0 u1 0 2.5463883302324e-06
Rx277 x277 0 1
Fxc277_278 x277 0 Vx278 767.385836045775
Cx277 x277 xm277 1.50857262477048e-14
Vx277 xm277 0 0
Gx277_1 x277 0 u1 0 -1.90876085584202e-09
Rx278 x278 0 1
Fxc278_277 x278 0 Vx277 -3451.20963066883
Cx278 x278 xm278 1.50857262477048e-14
Vx278 xm278 0 0
Gx278_1 x278 0 u1 0 6.58753384832567e-06
Rx279 x279 0 1
Fxc279_280 x279 0 Vx280 2960.49073293609
Cx279 x279 xm279 4.3895710802095e-15
Vx279 xm279 0 0
Gx279_1 x279 0 u1 0 -3.37910090863266e-10
Rx280 x280 0 1
Fxc280_279 x280 0 Vx279 -10628.6502640652
Cx280 x280 xm280 4.3895710802095e-15
Vx280 xm280 0 0
Gx280_1 x280 0 u1 0 3.59152817648414e-06
Rx281 x281 0 1
Fxc281_282 x281 0 Vx282 285.73331728064
Cx281 x281 xm281 1.55436740149653e-13
Vx281 xm281 0 0
Gx281_1 x281 0 u1 0 -2.03488763822199e-06
Rx282 x282 0 1
Fxc282_281 x282 0 Vx281 -89.2368983950997
Cx282 x282 xm282 1.55436740149653e-13
Vx282 xm282 0 0
Gx282_1 x282 0 u1 0 0.00018158706141746
Rx283 x283 0 1
Fxc283_284 x283 0 Vx284 8349.01574777647
Cx283 x283 xm283 1.56758610576001e-15
Vx283 xm283 0 0
Gx283_1 x283 0 u1 0 -3.95447313849019e-11
Rx284 x284 0 1
Fxc284_283 x284 0 Vx283 -29869.0982574649
Cx284 x284 xm284 1.56758610576001e-15
Vx284 xm284 0 0
Gx284_1 x284 0 u1 0 1.18116546730069e-06
Rx285 x285 0 1
Fxc285_286 x285 0 Vx286 84.4987875887279
Cx285 x285 xm285 3.97098834480777e-13
Vx285 xm285 0 0
Gx285_1 x285 0 u1 0 -4.79040432778738e-05
Rx286 x286 0 1
Fxc286_285 x286 0 Vx285 -48.0549950896333
Cx286 x286 xm286 3.97098834480777e-13
Vx286 xm286 0 0
Gx286_1 x286 0 u1 0 0.00230202856449181
Rx287 x287 0 1
Fxc287_288 x287 0 Vx288 33293.2782402952
Cx287 x287 xm287 1.20476536006176e-14
Vx287 xm287 0 0
Gx287_1 x287 0 u1 0 -5.89060383519489e-09
Rx288 x288 0 1
Fxc288_287 x288 0 Vx287 -127.583688119061
Cx288 x288 xm288 1.20476536006176e-14
Vx288 xm288 0 0
Gx288_1 x288 0 u1 0 7.51544962542447e-07
Rx289 x289 0 1
Fxc289_290 x289 0 Vx290 95066.3286437644
Cx289 x289 xm289 2.12416893515056e-16
Vx289 xm289 0 0
Gx289_1 x289 0 u1 0 -5.072512520865e-11
Rx290 x290 0 1
Fxc290_289 x290 0 Vx289 -146439.603232093
Cx290 x290 xm290 2.12416893515056e-16
Vx290 xm290 0 0
Gx290_1 x290 0 u1 0 7.42816720945295e-06
Rx291 x291 0 1
Fxc291_292 x291 0 Vx292 602.258228601248
Cx291 x291 xm291 9.7618575178155e-14
Vx291 xm291 0 0
Gx291_1 x291 0 u1 0 -5.41365282822917e-07
Rx292 x292 0 1
Fxc292_291 x292 0 Vx291 -109.784224512546
Cx292 x292 xm292 9.7618575178155e-14
Vx292 xm292 0 0
Gx292_1 x292 0 u1 0 5.9433367752729e-05
Rx293 x293 0 1
Fxc293_294 x293 0 Vx294 21202.4062699078
Cx293 x293 xm293 1.87292384452854e-15
Vx293 xm293 0 0
Gx293_1 x293 0 u1 0 -4.33472583856564e-10
Rx294 x294 0 1
Fxc294_293 x294 0 Vx293 -8604.89140864632
Cx294 x294 xm294 1.87292384452854e-15
Vx294 xm294 0 0
Gx294_1 x294 0 u1 0 3.72998451271107e-06
Rx295 x295 0 1
Fxc295_296 x295 0 Vx296 2053.32759132893
Cx295 x295 xm295 1.43078355234661e-14
Vx295 xm295 0 0
Gx295_1 x295 0 u1 0 -2.30216309805945e-08
Rx296 x296 0 1
Fxc296_295 x296 0 Vx295 -1522.4036857666
Cx296 x296 xm296 1.43078355234661e-14
Vx296 xm296 0 0
Gx296_1 x296 0 u1 0 3.50482158572155e-05
Rx297 x297 0 1
Fxc297_298 x297 0 Vx298 125.163132529755
Cx297 x297 xm297 1.25017605588615e-13
Vx297 xm297 0 0
Gx297_1 x297 0 u1 0 -8.69020056509006e-07
Rx298 x298 0 1
Fxc298_297 x298 0 Vx297 -369.566700522586
Cx298 x298 xm298 1.25017605588615e-13
Vx298 xm298 0 0
Gx298_1 x298 0 u1 0 0.000321160874971985
Rx299 x299 0 1
Fxc299_300 x299 0 Vx300 2024.53615745441
Cx299 x299 xm299 2.53678675984263e-14
Vx299 xm299 0 0
Gx299_1 x299 0 u1 0 -1.73093260488455e-08
Rx300 x300 0 1
Fxc300_299 x300 0 Vx299 -497.625941300819
Cx300 x300 xm300 2.53678675984263e-14
Vx300 xm300 0 0
Gx300_1 x300 0 u1 0 8.61356966833954e-06
Rx301 x301 0 1
Fxc301_302 x301 0 Vx302 166460.957957261
Cx301 x301 xm301 3.20804739778187e-16
Vx301 xm301 0 0
Gx301_1 x301 0 u1 0 -1.05704569199856e-10
Rx302 x302 0 1
Fxc302_301 x302 0 Vx301 -38017.737761674
Cx302 x302 xm302 3.20804739778187e-16
Vx302 xm302 0 0
Gx302_1 x302 0 u1 0 4.01864859205086e-06
Rx303 x303 0 1
Fxc303_304 x303 0 Vx304 12319.1097280921
Cx303 x303 xm303 2.27190048287476e-14
Vx303 xm303 0 0
Gx303_1 x303 0 u1 0 -1.00596767584225e-08
Rx304 x304 0 1
Fxc304_303 x304 0 Vx303 -103.490562291327
Cx304 x304 xm304 2.27190048287476e-14
Vx304 xm304 0 0
Gx304_1 x304 0 u1 0 1.04108160419814e-06
Rx305 x305 0 1
Fxc305_306 x305 0 Vx306 177.211132389894
Cx305 x305 xm305 2.2084230164543e-13
Vx305 xm305 0 0
Gx305_1 x305 0 u1 0 -8.69345516708659e-06
Rx306 x306 0 1
Fxc306_305 x306 0 Vx305 -78.346815453534
Cx306 x306 xm306 2.2084230164543e-13
Vx306 xm306 0 0
Gx306_1 x306 0 u1 0 0.000681104527629305
Rx307 x307 0 1
Fxc307_308 x307 0 Vx308 360.002800367105
Cx307 x307 xm307 2.43012562210102e-13
Vx307 xm307 0 0
Gx307_1 x307 0 u1 0 -1.16576239298203e-05
Rx308 x308 0 1
Fxc308_307 x308 0 Vx307 -32.5482132959345
Cx308 x308 xm308 2.43012562210102e-13
Vx308 xm308 0 0
Gx308_1 x308 0 u1 0 0.000379434830191582
Rx309 x309 0 1
Fxc309_310 x309 0 Vx310 1081.18783321622
Cx309 x309 xm309 3.92393390132605e-14
Vx309 xm309 0 0
Gx309_1 x309 0 u1 0 -3.64322563229217e-08
Rx310 x310 0 1
Fxc310_309 x310 0 Vx309 -406.533674452582
Cx310 x310 xm310 3.92393390132605e-14
Vx310 xm310 0 0
Gx310_1 x310 0 u1 0 1.48109390315557e-05
Rx311 x311 0 1
Fxc311_312 x311 0 Vx312 398.614470146252
Cx311 x311 xm311 2.14454644620413e-14
Vx311 xm311 0 0
Gx311_1 x311 0 u1 0 -3.55933029305661e-09
Rx312 x312 0 1
Fxc312_311 x312 0 Vx311 -3651.43714974526
Cx312 x312 xm312 2.14454644620413e-14
Vx312 xm312 0 0
Gx312_1 x312 0 u1 0 1.29966708602806e-05
Rx313 x313 0 1
Fxc313_314 x313 0 Vx314 33.9354038711674
Cx313 x313 xm313 3.69189637458766e-14
Vx313 xm313 0 0
Gx313_1 x313 0 u1 0 -1.70218412925843e-09
Rx314 x314 0 1
Fxc314_313 x314 0 Vx313 -14884.9140852841
Cx314 x314 xm314 3.69189637458766e-14
Vx314 xm314 0 0
Gx314_1 x314 0 u1 0 2.53368645213458e-05
Rx315 x315 0 1
Fxc315_316 x315 0 Vx316 1747.93011999887
Cx315 x315 xm315 1.78601578922452e-14
Vx315 xm315 0 0
Gx315_1 x315 0 u1 0 -4.83763175934404e-09
Rx316 x316 0 1
Fxc316_315 x316 0 Vx315 -1271.81933194008
Cx316 x316 xm316 1.78601578922452e-14
Vx316 xm316 0 0
Gx316_1 x316 0 u1 0 6.15259359234106e-06
Rx317 x317 0 1
Fxc317_318 x317 0 Vx318 6707.37133812251
Cx317 x317 xm317 3.02453155184689e-14
Vx317 xm317 0 0
Gx317_1 x317 0 u1 0 -1.83847498751122e-08
Rx318 x318 0 1
Fxc318_317 x318 0 Vx317 -113.183583693392
Cx318 x318 xm318 3.02453155184689e-14
Vx318 xm318 0 0
Gx318_1 x318 0 u1 0 2.08085187617185e-06
Rx319 x319 0 1
Fxc319_320 x319 0 Vx320 164.408610554148
Cx319 x319 xm319 3.68500092864944e-14
Vx319 xm319 0 0
Gx319_1 x319 0 u1 0 -5.81838478817977e-09
Rx320 x320 0 1
Fxc320_319 x320 0 Vx319 -3205.01341578256
Cx320 x320 xm320 3.68500092864944e-14
Vx320 xm320 0 0
Gx320_1 x320 0 u1 0 1.86480013043013e-05
Rx321 x321 0 1
Fxc321_322 x321 0 Vx322 660.789318115517
Cx321 x321 xm321 4.62675941996372e-14
Vx321 xm321 0 0
Gx321_1 x321 0 u1 0 -5.16559242850803e-08
Rx322 x322 0 1
Fxc322_321 x322 0 Vx321 -469.402859017121
Cx322 x322 xm322 4.62675941996372e-14
Vx322 xm322 0 0
Gx322_1 x322 0 u1 0 2.42474385445886e-05
Rx323 x323 0 1
Fxc323_324 x323 0 Vx324 7255.42414521675
Cx323 x323 xm323 2.94176684113735e-15
Vx323 xm323 0 0
Gx323_1 x323 0 u1 0 -3.07112980372767e-10
Rx324 x324 0 1
Fxc324_323 x324 0 Vx323 -11185.5161094648
Cx324 x324 xm324 2.94176684113735e-15
Vx324 xm324 0 0
Gx324_1 x324 0 u1 0 3.43521718938534e-06
Rx325 x325 0 1
Fxc325_326 x325 0 Vx326 1633.64220647998
Cx325 x325 xm325 9.26868572070505e-15
Vx325 xm325 0 0
Gx325_1 x325 0 u1 0 -1.60858861612801e-09
Rx326 x326 0 1
Fxc326_325 x326 0 Vx325 -5349.03648913451
Cx326 x326 xm326 9.26868572070505e-15
Vx326 xm326 0 0
Gx326_1 x326 0 u1 0 8.60439920367511e-06
Rx327 x327 0 1
Fxc327_328 x327 0 Vx328 674.67748317822
Cx327 x327 xm327 4.05009397042418e-14
Vx327 xm327 0 0
Gx327_1 x327 0 u1 0 -2.16101085611895e-08
Rx328 x328 0 1
Fxc328_327 x328 0 Vx327 -671.571769193826
Cx328 x328 xm328 4.05009397042418e-14
Vx328 xm328 0 0
Gx328_1 x328 0 u1 0 1.45127388389087e-05
Rx329 x329 0 1
Fxc329_330 x329 0 Vx330 10256.4194695901
Cx329 x329 xm329 4.03994326186591e-15
Vx329 xm329 0 0
Gx329_1 x329 0 u1 0 -7.32945014390107e-10
Rx330 x330 0 1
Fxc330_329 x330 0 Vx329 -4399.50789831542
Cx330 x330 xm330 4.03994326186591e-15
Vx330 xm330 0 0
Gx330_1 x330 0 u1 0 3.22459737984019e-06
Rx331 x331 0 1
Fxc331_332 x331 0 Vx332 4112.3945988542
Cx331 x331 xm331 1.4939511468885e-13
Vx331 xm331 0 0
Gx331_1 x331 0 u1 0 -3.03921398015573e-06
Rx332 x332 0 1
Fxc332_331 x332 0 Vx331 -7.91889951419369
Cx332 x332 xm332 1.4939511468885e-13
Vx332 xm332 0 0
Gx332_1 x332 0 u1 0 2.40672301109859e-05
Rx333 x333 0 1
Fxc333_334 x333 0 Vx334 4513.8707497803
Cx333 x333 xm333 1.24148427126151e-14
Vx333 xm333 0 0
Gx333_1 x333 0 u1 0 -2.18030575710432e-09
Rx334 x334 0 1
Fxc334_333 x334 0 Vx333 -1043.48866491322
Cx334 x334 xm334 1.24148427126151e-14
Vx334 xm334 0 0
Gx334_1 x334 0 u1 0 2.2751243435834e-06
Rx335 x335 0 1
Fxc335_336 x335 0 Vx336 926.515322261138
Cx335 x335 xm335 3.04285853351407e-14
Vx335 xm335 0 0
Gx335_1 x335 0 u1 0 -1.21719533276507e-08
Rx336 x336 0 1
Fxc336_335 x336 0 Vx335 -884.194447463008
Cx336 x336 xm336 3.04285853351407e-14
Vx336 xm336 0 0
Gx336_1 x336 0 u1 0 1.07623735470876e-05
Rx337 x337 0 1
Fxc337_338 x337 0 Vx338 82886.1112909633
Cx337 x337 xm337 2.80028892882111e-16
Vx337 xm337 0 0
Gx337_1 x337 0 u1 0 -1.43225612376604e-11
Rx338 x338 0 1
Fxc338_337 x338 0 Vx337 -118297.892621305
Cx338 x338 xm338 2.80028892882111e-16
Vx338 xm338 0 0
Gx338_1 x338 0 u1 0 1.69432881135482e-06
Rx339 x339 0 1
Fxc339_340 x339 0 Vx340 7318.16663819316
Cx339 x339 xm339 5.53119643557016e-15
Vx339 xm339 0 0
Gx339_1 x339 0 u1 0 -7.456270034575e-10
Rx340 x340 0 1
Fxc340_339 x340 0 Vx339 -3504.1172226728
Cx340 x340 xm340 5.53119643557016e-15
Vx340 xm340 0 0
Gx340_1 x340 0 u1 0 2.61276442450534e-06
Rx341 x341 0 1
Fxc341_342 x341 0 Vx342 22263.1460632585
Cx341 x341 xm341 3.62906157244733e-15
Vx341 xm341 0 0
Gx341_1 x341 0 u1 0 -3.38067382020427e-10
Rx342 x342 0 1
Fxc342_341 x342 0 Vx341 -2646.41599476803
Cx342 x342 xm342 3.62906157244733e-15
Vx342 xm342 0 0
Gx342_1 x342 0 u1 0 8.94666927088211e-07
Rx343 x343 0 1
Fxc343_344 x343 0 Vx344 1307.42825718444
Cx343 x343 xm343 2.43563137386751e-14
Vx343 xm343 0 0
Gx343_1 x343 0 u1 0 -7.4034295004626e-09
Rx344 x344 0 1
Fxc344_343 x344 0 Vx343 -1027.81849331455
Cx344 x344 xm344 2.43563137386751e-14
Vx344 xm344 0 0
Gx344_1 x344 0 u1 0 7.60938175452596e-06
Rx345 x345 0 1
Fxc345_346 x345 0 Vx346 11853.1271774998
Cx345 x345 xm345 7.64511008833616e-15
Vx345 xm345 0 0
Gx345_1 x345 0 u1 0 -6.92845986252749e-10
Rx346 x346 0 1
Fxc346_345 x346 0 Vx345 -1143.77278805996
Cx346 x346 xm346 7.64511008833616e-15
Vx346 xm346 0 0
Gx346_1 x346 0 u1 0 7.92458385392459e-07
Rx347 x347 0 1
Fxc347_348 x347 0 Vx348 263.651585569789
Cx347 x347 xm347 3.31932360252982e-14
Vx347 xm347 0 0
Gx347_1 x347 0 u1 0 -8.25858693325056e-09
Rx348 x348 0 1
Fxc348_347 x348 0 Vx347 -2599.9044126119
Cx348 x348 xm348 3.31932360252982e-14
Vx348 xm348 0 0
Gx348_1 x348 0 u1 0 2.14715366096971e-05
Rx349 x349 0 1
Fxc349_350 x349 0 Vx350 52.0283492581108
Cx349 x349 xm349 3.91990471759038e-13
Vx349 xm349 0 0
Gx349_1 x349 0 u1 0 -5.12033316777386e-05
Rx350 x350 0 1
Fxc350_349 x350 0 Vx349 -103.887553155089
Cx350 x350 xm350 3.91990471759038e-13
Vx350 xm350 0 0
Gx350_1 x350 0 u1 0 0.00531938884138871
Rx351 x351 0 1
Fxc351_352 x351 0 Vx352 3802.73051282273
Cx351 x351 xm351 1.62720964829041e-14
Vx351 xm351 0 0
Gx351_1 x351 0 u1 0 -9.02205122199579e-09
Rx352 x352 0 1
Fxc352_351 x352 0 Vx351 -799.675739241955
Cx352 x352 xm352 1.62720964829041e-14
Vx352 xm352 0 0
Gx352_1 x352 0 u1 0 7.21471548042827e-06
Rx353 x353 0 1
Fxc353_354 x353 0 Vx354 3616.65361389252
Cx353 x353 xm353 8.80522494224566e-14
Vx353 xm353 0 0
Gx353_1 x353 0 u1 0 -3.49502620448498e-07
Rx354 x354 0 1
Fxc354_353 x354 0 Vx353 -28.7367320045547
Cx354 x354 xm354 8.80522494224566e-14
Vx354 xm354 0 0
Gx354_1 x354 0 u1 0 1.00435631387181e-05
Rx355 x355 0 1
Fxc355_356 x355 0 Vx356 7.12868110480384
Cx355 x355 xm355 7.67229662280685e-13
Vx355 xm355 0 0
Gx355_1 x355 0 u1 0 -0.000100857350424888
Rx356 x356 0 1
Fxc356_355 x356 0 Vx355 -214.691370393248
Cx356 x356 xm356 7.67229662280685e-13
Vx356 xm356 0 0
Gx356_1 x356 0 u1 0 0.0216532027769512
Rx357 x357 0 1
Fxc357_358 x357 0 Vx358 8.55688336515506
Cx357 x357 xm357 4.92776735733474e-13
Vx357 xm357 0 0
Gx357_1 x357 0 u1 0 -3.13220807637156e-05
Rx358 x358 0 1
Fxc358_357 x358 0 Vx357 -402.347204487387
Cx358 x358 xm358 4.92776735733474e-13
Vx358 xm358 0 0
Gx358_1 x358 0 u1 0 0.0126023516340091
Rx359 x359 0 1
Fxc359_360 x359 0 Vx360 1406.72586024309
Cx359 x359 xm359 1.65994637491899e-14
Vx359 xm359 0 0
Gx359_1 x359 0 u1 0 -1.90154325241204e-09
Rx360 x360 0 1
Fxc360_359 x360 0 Vx359 -2110.22251723069
Cx360 x360 xm360 1.65994637491899e-14
Vx360 xm360 0 0
Gx360_1 x360 0 u1 0 4.01267938872796e-06
Rx361 x361 0 1
Fxc361_362 x361 0 Vx362 333.49377827196
Cx361 x361 xm361 1.52443737477815e-14
Vx361 xm361 0 0
Gx361_1 x361 0 u1 0 -1.4040109440449e-10
Rx362 x362 0 1
Fxc362_361 x362 0 Vx361 -10650.5648089138
Cx362 x362 xm362 1.52443737477815e-14
Vx362 xm362 0 0
Gx362_1 x362 0 u1 0 1.49535095519745e-06
Rx363 x363 0 1
Fxc363_364 x363 0 Vx364 114.73896077935
Cx363 x363 xm363 2.73296090832205e-13
Vx363 xm363 0 0
Gx363_1 x363 0 u1 0 -9.93421377831721e-06
Rx364 x364 0 1
Fxc364_363 x364 0 Vx363 -106.956620327395
Cx364 x364 xm364 2.73296090832205e-13
Vx364 xm364 0 0
Gx364_1 x364 0 u1 0 0.00106252993133865
Rx365 x365 0 1
Fxc365_366 x365 0 Vx366 737.879180772056
Cx365 x365 xm365 2.87228473774017e-14
Vx365 xm365 0 0
Gx365_1 x365 0 u1 0 -5.69552654953577e-09
Rx366 x366 0 1
Fxc366_365 x366 0 Vx365 -1380.33774930498
Cx366 x366 xm366 2.87228473774017e-14
Vx366 xm366 0 0
Gx366_1 x366 0 u1 0 7.86175029849296e-06
Rx367 x367 0 1
Fxc367_368 x367 0 Vx368 1102.13015435471
Cx367 x367 xm367 4.66685567425351e-14
Vx367 xm367 0 0
Gx367_1 x367 0 u1 0 -3.61427415383075e-08
Rx368 x368 0 1
Fxc368_367 x368 0 Vx367 -354.883160915616
Cx368 x368 xm368 4.66685567425351e-14
Vx368 xm368 0 0
Gx368_1 x368 0 u1 0 1.28264503612707e-05
Rx369 x369 0 1
Fxc369_370 x369 0 Vx370 949.658661832279
Cx369 x369 xm369 5.7196013910315e-14
Vx369 xm369 0 0
Gx369_1 x369 0 u1 0 -6.98854487157505e-08
Rx370 x370 0 1
Fxc370_369 x370 0 Vx369 -276.34279737955
Cx370 x370 xm370 5.7196013910315e-14
Vx370 xm370 0 0
Gx370_1 x370 0 u1 0 1.93123403942356e-05
Rx371 x371 0 1
Fxc371_372 x371 0 Vx372 230.947965874743
Cx371 x371 xm371 1.75688323351063e-13
Vx371 xm371 0 0
Gx371_1 x371 0 u1 0 -2.85150700570423e-06
Rx372 x372 0 1
Fxc372_371 x372 0 Vx371 -124.428064768907
Cx372 x372 xm372 1.75688323351063e-13
Vx372 xm372 0 0
Gx372_1 x372 0 u1 0 0.000354807498394757
Rx373 x373 0 1
Fxc373_374 x373 0 Vx374 13124.4601806389
Cx373 x373 xm373 6.22004467114814e-14
Vx373 xm373 0 0
Gx373_1 x373 0 u1 0 -9.62578860956846e-08
Rx374 x374 0 1
Fxc374_373 x374 0 Vx373 -17.62577564018
Cx374 x374 xm374 6.22004467114814e-14
Vx374 xm374 0 0
Gx374_1 x374 0 u1 0 1.69661990392054e-06
Rx375 x375 0 1
Fxc375_376 x375 0 Vx376 5627.54474829777
Cx375 x375 xm375 1.41434995567386e-14
Vx375 xm375 0 0
Gx375_1 x375 0 u1 0 -2.43423907290962e-09
Rx376 x376 0 1
Fxc376_375 x376 0 Vx375 -774.074571810792
Cx376 x376 xm376 1.41434995567386e-14
Vx376 xm376 0 0
Gx376_1 x376 0 u1 0 1.88428256804761e-06
Rx377 x377 0 1
Fxc377_378 x377 0 Vx378 257.39448937113
Cx377 x377 xm377 5.26768043602151e-14
Vx377 xm377 0 0
Gx377_1 x377 0 u1 0 -2.61484416046451e-08
Rx378 x378 0 1
Fxc378_377 x378 0 Vx377 -1233.67630057658
Cx378 x378 xm378 5.26768043602151e-14
Vx378 xm378 0 0
Gx378_1 x378 0 u1 0 3.22587127046614e-05
Rx379 x379 0 1
Fxc379_380 x379 0 Vx380 1482.91831880754
Cx379 x379 xm379 5.31047753536345e-14
Vx379 xm379 0 0
Gx379_1 x379 0 u1 0 -4.5934958461747e-08
Rx380 x380 0 1
Fxc380_379 x380 0 Vx379 -217.564296261868
Cx380 x380 xm380 5.31047753536345e-14
Vx380 xm380 0 0
Gx380_1 x380 0 u1 0 9.99380691154813e-06
Rx381 x381 0 1
Fxc381_382 x381 0 Vx382 1062.96653553824
Cx381 x381 xm381 1.32036835764334e-14
Vx381 xm381 0 0
Gx381_1 x381 0 u1 0 -2.74622328593114e-10
Rx382 x382 0 1
Fxc382_381 x382 0 Vx381 -4968.0706645205
Cx382 x382 xm382 1.32036835764334e-14
Vx382 xm382 0 0
Gx382_1 x382 0 u1 0 1.36434313450576e-06
Rx383 x383 0 1
Fxc383_384 x383 0 Vx384 36.3002173548474
Cx383 x383 xm383 5.7822019650203e-13
Vx383 xm383 0 0
Gx383_1 x383 0 u1 0 -0.000114182603522677
Rx384 x384 0 1
Fxc384_383 x384 0 Vx383 -80.8152531310451
Cx384 x384 xm384 5.7822019650203e-13
Vx384 xm384 0 0
Gx384_1 x384 0 u1 0 0.0092276960068469
Rx385 x385 0 1
Fxc385_386 x385 0 Vx386 563.482268777598
Cx385 x385 xm385 1.02035760349352e-13
Vx385 xm385 0 0
Gx385_1 x385 0 u1 0 -3.40428655145676e-07
Rx386 x386 0 1
Fxc386_385 x386 0 Vx385 -159.025939604156
Cx386 x386 xm386 1.02035760349352e-13
Vx386 xm386 0 0
Gx386_1 x386 0 u1 0 5.41369867527204e-05
Rx387 x387 0 1
Fxc387_388 x387 0 Vx388 3649.51279750134
Cx387 x387 xm387 2.40247346728811e-14
Vx387 xm387 0 0
Gx387_1 x387 0 u1 0 -1.03479335299402e-08
Rx388 x388 0 1
Fxc388_387 x388 0 Vx387 -447.354604662377
Cx388 x388 xm388 2.40247346728811e-14
Vx388 xm388 0 0
Gx388_1 x388 0 u1 0 4.62919571335897e-06
Rx389 x389 0 1
Fxc389_390 x389 0 Vx390 144.110234409434
Cx389 x389 xm389 3.08852421707331e-14
Vx389 xm389 0 0
Gx389_1 x389 0 u1 0 -1.46826134511536e-09
Rx390 x390 0 1
Fxc390_389 x390 0 Vx389 -6920.93971884088
Cx390 x390 xm390 3.08852421707331e-14
Vx390 xm390 0 0
Gx390_1 x390 0 u1 0 1.01617482610476e-05
Rx391 x391 0 1
Fxc391_392 x391 0 Vx392 477.922545101204
Cx391 x391 xm391 1.63019845419542e-14
Vx391 xm391 0 0
Gx391_1 x391 0 u1 0 -7.18725977975989e-10
Rx392 x392 0 1
Fxc392_391 x392 0 Vx391 -7541.14895133774
Cx392 x392 xm392 1.63019845419542e-14
Vx392 xm392 0 0
Gx392_1 x392 0 u1 0 5.42001965511281e-06
Rx393 x393 0 1
Fxc393_394 x393 0 Vx394 97.0221149376874
Cx393 x393 xm393 6.41736383827721e-13
Vx393 xm393 0 0
Gx393_1 x393 0 u1 0 -0.000168422901227077
Rx394 x394 0 1
Fxc394_393 x394 0 Vx393 -26.251838875632
Cx394 x394 xm394 6.41736383827721e-13
Vx394 xm394 0 0
Gx394_1 x394 0 u1 0 0.0044214108659797
Rx395 x395 0 1
Fxc395_396 x395 0 Vx396 184.359478877959
Cx395 x395 xm395 2.85479875469681e-14
Vx395 xm395 0 0
Gx395_1 x395 0 u1 0 -1.79648017094755e-09
Rx396 x396 0 1
Fxc396_395 x396 0 Vx395 -6451.17676952365
Cx396 x396 xm396 2.85479875469681e-14
Vx396 xm396 0 0
Gx396_1 x396 0 u1 0 1.15894111457267e-05
Rx397 x397 0 1
Fxc397_398 x397 0 Vx398 28.7592824344018
Cx397 x397 xm397 5.3285703820123e-13
Vx397 xm397 0 0
Gx397_1 x397 0 u1 0 -9.23163600772872e-05
Rx398 x398 0 1
Fxc398_397 x398 0 Vx397 -123.903741533266
Cx398 x398 xm398 5.3285703820123e-13
Vx398 xm398 0 0
Gx398_1 x398 0 u1 0 0.0114383424183081
Rx399 x399 0 1
Fxc399_400 x399 0 Vx400 203.581322180354
Cx399 x399 xm399 3.03498701128083e-14
Vx399 xm399 0 0
Gx399_1 x399 0 u1 0 -2.15015241680905e-09
Rx400 x400 0 1
Fxc400_399 x400 0 Vx399 -5201.77884695275
Cx400 x400 xm400 3.03498701128083e-14
Vx400 xm400 0 0
Gx400_1 x400 0 u1 0 1.11846173594817e-05
Rx401 x401 0 1
Fxc401_402 x401 0 Vx402 488.90943112262
Cx401 x401 xm401 1.01462685758652e-13
Vx401 xm401 0 0
Gx401_1 x401 0 u1 0 -3.19940714635596e-07
Rx402 x402 0 1
Fxc402_401 x402 0 Vx401 -197.908410345252
Cx402 x402 xm402 1.01462685758652e-13
Vx402 xm402 0 0
Gx402_1 x402 0 u1 0 6.33189582382549e-05
Rx403 x403 0 1
Fxc403_404 x403 0 Vx404 1156.38389683199
Cx403 x403 xm403 1.02325988713972e-13
Vx403 xm403 0 0
Gx403_1 x403 0 u1 0 -3.97232529812939e-07
Rx404 x404 0 1
Fxc404_403 x404 0 Vx403 -83.0894934071482
Cx404 x404 xm404 1.02325988713972e-13
Vx404 xm404 0 0
Gx404_1 x404 0 u1 0 3.3005849666997e-05
Rx405 x405 0 1
Fxc405_406 x405 0 Vx406 125.269816106537
Cx405 x405 xm405 1.41000112840634e-13
Vx405 xm405 0 0
Gx405_1 x405 0 u1 0 -1.39484580251953e-06
Rx406 x406 0 1
Fxc406_405 x406 0 Vx405 -457.318416400801
Cx406 x406 xm406 1.41000112840634e-13
Vx406 xm406 0 0
Gx406_1 x406 0 u1 0 0.000637888673531538
Rx407 x407 0 1
Fxc407_408 x407 0 Vx408 241.752050967692
Cx407 x407 xm407 1.32754836741219e-13
Vx407 xm407 0 0
Gx407_1 x407 0 u1 0 -4.37061535893652e-07
Rx408 x408 0 1
Fxc408_407 x408 0 Vx407 -240.449673699553
Cx408 x408 xm408 1.32754836741219e-13
Vx408 xm408 0 0
Gx408_1 x408 0 u1 0 0.000105091303692254
Rx409 x409 0 1
Fxc409_410 x409 0 Vx410 2676.84481459112
Cx409 x409 xm409 1.26702180135926e-14
Vx409 xm409 0 0
Gx409_1 x409 0 u1 0 -2.41901838638444e-09
Rx410 x410 0 1
Fxc410_409 x410 0 Vx409 -2615.05593595835
Cx410 x410 xm410 1.26702180135926e-14
Vx410 xm410 0 0
Gx410_1 x410 0 u1 0 6.32586839050701e-06
Rx411 x411 0 1
Fxc411_412 x411 0 Vx412 129.707208429803
Cx411 x411 xm411 3.01789464736231e-14
Vx411 xm411 0 0
Gx411_1 x411 0 u1 0 -9.86442829507094e-10
Rx412 x412 0 1
Fxc412_411 x412 0 Vx411 -8992.69222213537
Cx412 x412 xm412 3.01789464736231e-14
Vx412 xm412 0 0
Gx412_1 x412 0 u1 0 8.87077676048965e-06
Rx413 x413 0 1
Fxc413_414 x413 0 Vx414 1266.08340007649
Cx413 x413 xm413 9.70484385291883e-14
Vx413 xm413 0 0
Gx413_1 x413 0 u1 0 -5.06879481039693e-07
Rx414 x414 0 1
Fxc414_413 x414 0 Vx413 -91.7922830566829
Cx414 x414 xm414 9.70484385291882e-14
Vx414 xm414 0 0
Gx414_1 x414 0 u1 0 4.652762479922e-05
Rx415 x415 0 1
Fxc415_416 x415 0 Vx416 825.649940955848
Cx415 x415 xm415 3.43607207471199e-14
Vx415 xm415 0 0
Gx415_1 x415 0 u1 0 -9.69616718015153e-09
Rx416 x416 0 1
Fxc416_415 x416 0 Vx415 -1082.18045256972
Cx416 x416 xm416 3.43607207471199e-14
Vx416 xm416 0 0
Gx416_1 x416 0 u1 0 1.0493002587208e-05
Rx417 x417 0 1
Fxc417_418 x417 0 Vx418 241.665773765583
Cx417 x417 xm417 1.54871227469822e-13
Vx417 xm417 0 0
Gx417_1 x417 0 u1 0 -1.72883842020163e-06
Rx418 x418 0 1
Fxc418_417 x418 0 Vx417 -189.801075515044
Cx418 x418 xm418 1.54871227469822e-13
Vx418 xm418 0 0
Gx418_1 x418 0 u1 0 0.000328135391545999
Rx419 x419 0 1
Fxc419_420 x419 0 Vx420 39.1682572162851
Cx419 x419 xm419 6.44307967443506e-14
Vx419 xm419 0 0
Gx419_1 x419 0 u1 0 -4.2798008162292e-09
Rx420 x420 0 1
Fxc420_419 x420 0 Vx419 -6654.51521178315
Cx420 x420 xm420 6.44307967443506e-14
Vx420 xm420 0 0
Gx420_1 x420 0 u1 0 2.84799996349992e-05
Rx421 x421 0 1
Fxc421_422 x421 0 Vx422 5529.41673512099
Cx421 x421 xm421 2.24357038343354e-14
Vx421 xm421 0 0
Gx421_1 x421 0 u1 0 -1.56050339748984e-08
Rx422 x422 0 1
Fxc422_421 x422 0 Vx421 -394.874214610616
Cx422 x422 xm422 2.24357038343354e-14
Vx422 xm422 0 0
Gx422_1 x422 0 u1 0 6.16202553481001e-06
Rx423 x423 0 1
Fxc423_424 x423 0 Vx424 84.9086267080667
Cx423 x423 xm423 2.99137106960636e-14
Vx423 xm423 0 0
Gx423_1 x423 0 u1 0 -3.99461027425459e-10
Rx424 x424 0 1
Fxc424_423 x424 0 Vx423 -13668.1401564053
Cx424 x424 xm424 2.99137106960636e-14
Vx424 xm424 0 0
Gx424_1 x424 0 u1 0 5.45988930987284e-06
Rx425 x425 0 1
Fxc425_426 x425 0 Vx426 107.509932367549
Cx425 x425 xm425 2.79263378446224e-13
Vx425 xm425 0 0
Gx425_1 x425 0 u1 0 -8.80087707283007e-06
Rx426 x426 0 1
Fxc426_425 x426 0 Vx425 -138.41645921036
Cx426 x426 xm426 2.79263378446224e-13
Vx426 xm426 0 0
Gx426_1 x426 0 u1 0 0.00121818624236677
Rx427 x427 0 1
Fxc427_428 x427 0 Vx428 185.255921124301
Cx427 x427 xm427 1.23092401377661e-13
Vx427 xm427 0 0
Gx427_1 x427 0 u1 0 -1.18808438328085e-06
Rx428 x428 0 1
Fxc428_427 x428 0 Vx427 -407.235383214653
Cx428 x428 xm428 1.23092401377661e-13
Vx428 xm428 0 0
Gx428_1 x428 0 u1 0 0.000483829999116721
Rx429 x429 0 1
Fxc429_430 x429 0 Vx430 4.60177108819814
Cx429 x429 xm429 2.82424764335851e-12
Vx429 xm429 0 0
Gx429_1 x429 0 u1 0 -0.00222597507611063
Rx430 x430 0 1
Fxc430_429 x430 0 Vx429 -35.426814276598
Cx430 x430 xm430 2.82424764335851e-12
Vx430 xm430 0 0
Gx430_1 x430 0 u1 0 0.0788592056057075
Rx431 x431 0 1
Fxc431_432 x431 0 Vx432 1029.33524139771
Cx431 x431 xm431 1.22590423162195e-13
Vx431 xm431 0 0
Gx431_1 x431 0 u1 0 -7.20426490713617e-07
Rx432 x432 0 1
Fxc432_431 x432 0 Vx431 -79.4105995904914
Cx432 x432 xm432 1.22590423162195e-13
Vx432 xm432 0 0
Gx432_1 x432 0 u1 0 5.72094995884419e-05
Rx433 x433 0 1
Fxc433_434 x433 0 Vx434 196.162743926585
Cx433 x433 xm433 4.09020191567389e-13
Vx433 xm433 0 0
Gx433_1 x433 0 u1 0 -3.35648464132663e-05
Rx434 x434 0 1
Fxc434_433 x434 0 Vx433 -37.2438898038179
Cx434 x434 xm434 4.09020191567389e-13
Vx434 xm434 0 0
Gx434_1 x434 0 u1 0 0.00125008544109776
Rx435 x435 0 1
Fxc435_436 x435 0 Vx436 5115.72026495366
Cx435 x435 xm435 9.93705359088137e-14
Vx435 xm435 0 0
Gx435_1 x435 0 u1 0 -5.07181960793568e-07
Rx436 x436 0 1
Fxc436_435 x436 0 Vx435 -23.8433646305929
Cx436 x436 xm436 9.93705359088137e-14
Vx436 xm436 0 0
Gx436_1 x436 0 u1 0 1.20929244252601e-05
Rx437 x437 0 1
Fxc437_438 x437 0 Vx438 311.300979434606
Cx437 x437 xm437 5.79622437737296e-14
Vx437 xm437 0 0
Gx437_1 x437 0 u1 0 -4.20297355468863e-08
Rx438 x438 0 1
Fxc438_437 x438 0 Vx437 -1110.36847871201
Cx438 x438 xm438 5.79622437737296e-14
Vx438 xm438 0 0
Gx438_1 x438 0 u1 0 4.66684935198642e-05
Rx439 x439 0 1
Fxc439_440 x439 0 Vx440 2286.41298552075
Cx439 x439 xm439 3.54576514760153e-14
Vx439 xm439 0 0
Gx439_1 x439 0 u1 0 -1.84228410539917e-08
Rx440 x440 0 1
Fxc440_439 x440 0 Vx439 -411.258666205796
Cx440 x440 xm440 3.54576514760153e-14
Vx440 xm440 0 0
Gx440_1 x440 0 u1 0 7.57655303958602e-06
Rx441 x441 0 1
Fxc441_442 x441 0 Vx442 147.183246513882
Cx441 x441 xm441 1.2896763528379e-13
Vx441 xm441 0 0
Gx441_1 x441 0 u1 0 -5.38636051905471e-07
Rx442 x442 0 1
Fxc442_441 x442 0 Vx441 -489.102057110588
Cx442 x442 xm442 1.2896763528379e-13
Vx442 xm442 0 0
Gx442_1 x442 0 u1 0 0.000263448001020891
Rx443 x443 0 1
Fxc443_444 x443 0 Vx444 941.902583479155
Cx443 x443 xm443 9.26424551985641e-14
Vx443 xm443 0 0
Gx443_1 x443 0 u1 0 -2.55054794845631e-07
Rx444 x444 0 1
Fxc444_443 x444 0 Vx443 -153.551520443144
Cx444 x444 xm444 9.26424551985641e-14
Vx444 xm444 0 0
Gx444_1 x444 0 u1 0 3.91640515448609e-05
Rx445 x445 0 1
Fxc445_446 x445 0 Vx446 5790.92767874224
Cx445 x445 xm445 1.72944646712239e-14
Vx445 xm445 0 0
Gx445_1 x445 0 u1 0 -4.17445562243291e-09
Rx446 x446 0 1
Fxc446_445 x446 0 Vx445 -723.478969051808
Cx446 x446 xm446 1.72944646712239e-14
Vx446 xm446 0 0
Gx446_1 x446 0 u1 0 3.02013085007029e-06
Rx447 x447 0 1
Fxc447_448 x447 0 Vx448 41.8033490863968
Cx447 x447 xm447 3.11153675188471e-13
Vx447 xm447 0 0
Gx447_1 x447 0 u1 0 -1.60855908927776e-06
Rx448 x448 0 1
Fxc448_447 x448 0 Vx447 -345.394856738367
Cx448 x448 xm448 3.11153675188471e-13
Vx448 xm448 0 0
Gx448_1 x448 0 u1 0 0.000555588036196289
Rx449 x449 0 1
Fxc449_450 x449 0 Vx450 69.4452698268554
Cx449 x449 xm449 4.37725075845039e-13
Vx449 xm449 0 0
Gx449_1 x449 0 u1 0 -1.28385019831166e-05
Rx450 x450 0 1
Fxc450_449 x450 0 Vx449 -102.849621768964
Cx450 x450 xm450 4.37725075845039e-13
Vx450 xm450 0 0
Gx450_1 x450 0 u1 0 0.00132043507304364
Rx451 x451 0 1
Fxc451_452 x451 0 Vx452 602.804567288196
Cx451 x451 xm451 2.89789505961041e-14
Vx451 xm451 0 0
Gx451_1 x451 0 u1 0 -4.49371230132991e-09
Rx452 x452 0 1
Fxc452_451 x452 0 Vx451 -2526.82778614825
Cx452 x452 xm452 2.89789505961041e-14
Vx452 xm452 0 0
Gx452_1 x452 0 u1 0 1.13548371059566e-05
Rx453 x453 0 1
Fxc453_454 x453 0 Vx454 35.5267146741572
Cx453 x453 xm453 3.08257267736937e-13
Vx453 xm453 0 0
Gx453_1 x453 0 u1 0 -1.88423756066304e-06
Rx454 x454 0 1
Fxc454_453 x454 0 Vx453 -390.176140184932
Cx454 x454 xm454 3.08257267736937e-13
Vx454 xm454 0 0
Gx454_1 x454 0 u1 0 0.000735184538610977
Rx455 x455 0 1
Fxc455_456 x455 0 Vx456 22035.7832480319
Cx455 x455 xm455 6.93829485175084e-14
Vx455 xm455 0 0
Gx455_1 x455 0 u1 0 -6.9784398515398e-08
Rx456 x456 0 1
Fxc456_455 x456 0 Vx455 -12.2272829126758
Cx456 x456 xm456 6.93829485175084e-14
Vx456 xm456 0 0
Gx456_1 x456 0 u1 0 8.53273583538686e-07
Rx457 x457 0 1
Fxc457_458 x457 0 Vx458 10.3561514542354
Cx457 x457 xm457 8.93653863244677e-14
Vx457 xm457 0 0
Gx457_1 x457 0 u1 0 -3.43893446970616e-09
Rx458 x458 0 1
Fxc458_457 x458 0 Vx457 -16451.9234242339
Cx458 x458 xm458 8.93653863244677e-14
Vx458 xm458 0 0
Gx458_1 x458 0 u1 0 5.65770865565643e-05
Rx459 x459 0 1
Fxc459_460 x459 0 Vx460 1307.18769053511
Cx459 x459 xm459 7.05517351858277e-14
Vx459 xm459 0 0
Gx459_1 x459 0 u1 0 -7.68709221587628e-08
Rx460 x460 0 1
Fxc460_459 x460 0 Vx459 -201.13014457431
Cx460 x460 xm460 7.05517351858277e-14
Vx460 xm460 0 0
Gx460_1 x460 0 u1 0 1.54610596873525e-05
Rx461 x461 0 1
Fxc461_462 x461 0 Vx462 517.849273745909
Cx461 x461 xm461 1.82509464382829e-14
Vx461 xm461 0 0
Gx461_1 x461 0 u1 0 -6.95414401646122e-10
Rx462 x462 0 1
Fxc462_461 x462 0 Vx461 -7970.67417935588
Cx462 x462 xm462 1.82509464382829e-14
Vx462 xm462 0 0
Gx462_1 x462 0 u1 0 5.54292161515296e-06
Rx463 x463 0 1
Fxc463_464 x463 0 Vx464 8771.14794482321
Cx463 x463 xm463 2.53969224170102e-14
Vx463 xm463 0 0
Gx463_1 x463 0 u1 0 -8.53613950787934e-09
Rx464 x464 0 1
Fxc464_463 x464 0 Vx463 -235.055438035171
Cx464 x464 xm464 2.53969224170102e-14
Vx464 xm464 0 0
Gx464_1 x464 0 u1 0 2.00646601115391e-06
Rx465 x465 0 1
Fxc465_466 x465 0 Vx466 9044.08719708216
Cx465 x465 xm465 2.15604352286956e-14
Vx465 xm465 0 0
Gx465_1 x465 0 u1 0 -8.7672826353503e-09
Rx466 x466 0 1
Fxc466_465 x466 0 Vx465 -335.270592650388
Cx466 x466 xm466 2.15604352286955e-14
Vx466 xm466 0 0
Gx466_1 x466 0 u1 0 2.93941204508735e-06
Rx467 x467 0 1
Fxc467_468 x467 0 Vx468 77.2231923138224
Cx467 x467 xm467 6.88076389610427e-14
Vx467 xm467 0 0
Gx467_1 x467 0 u1 0 -6.66072322270681e-09
Rx468 x468 0 1
Fxc468_467 x468 0 Vx467 -3908.81057929838
Cx468 x468 xm468 6.88076389610427e-14
Vx468 xm468 0 0
Gx468_1 x468 0 u1 0 2.60355053986948e-05
Rx469 x469 0 1
Fxc469_470 x469 0 Vx470 141.827713278729
Cx469 x469 xm469 3.36224705594798e-14
Vx469 xm469 0 0
Gx469_1 x469 0 u1 0 -1.57941340528927e-09
Rx470 x470 0 1
Fxc470_469 x470 0 Vx469 -9022.17932015636
Cx470 x470 xm470 3.36224705594798e-14
Vx470 xm470 0 0
Gx470_1 x470 0 u1 0 1.42497509631786e-05
Rx471 x471 0 1
Fxc471_472 x471 0 Vx472 1040.25567577254
Cx471 x471 xm471 3.82271448805577e-14
Vx471 xm471 0 0
Gx471_1 x471 0 u1 0 -7.45439376911983e-09
Rx472 x472 0 1
Fxc472_471 x472 0 Vx471 -970.675523578247
Cx472 x472 xm472 3.82271448805577e-14
Vx472 xm472 0 0
Gx472_1 x472 0 u1 0 7.23579757479882e-06
Rx473 x473 0 1
Fxc473_474 x473 0 Vx474 42.4555010312021
Cx473 x473 xm473 1.20061702453183e-13
Vx473 xm473 0 0
Gx473_1 x473 0 u1 0 -3.18645815322136e-08
Rx474 x474 0 1
Fxc474_473 x474 0 Vx473 -2462.11596342576
Cx474 x474 xm474 1.20061702453183e-13
Vx474 xm474 0 0
Gx474_1 x474 0 u1 0 7.84542948583446e-05
Rx475 x475 0 1
Fxc475_476 x475 0 Vx476 1290.33251720867
Cx475 x475 xm475 5.54932867986001e-14
Vx475 xm475 0 0
Gx475_1 x475 0 u1 0 -3.16950758397224e-08
Rx476 x476 0 1
Fxc476_475 x476 0 Vx475 -376.744029445715
Cx476 x476 xm476 5.54932867986001e-14
Vx476 xm476 0 0
Gx476_1 x476 0 u1 0 1.19409305854446e-05
Rx477 x477 0 1
Fxc477_478 x477 0 Vx478 170.633770669981
Cx477 x477 xm477 6.24009086699585e-14
Vx477 xm477 0 0
Gx477_1 x477 0 u1 0 -1.4908695196481e-08
Rx478 x478 0 1
Fxc478_477 x478 0 Vx477 -2293.23426023551
Cx478 x478 xm478 6.24009086699586e-14
Vx478 xm478 0 0
Gx478_1 x478 0 u1 0 3.41891305999787e-05
Rx479 x479 0 1
Fxc479_480 x479 0 Vx480 296.187270917459
Cx479 x479 xm479 6.64567064981729e-14
Vx479 xm479 0 0
Gx479_1 x479 0 u1 0 -2.87849984836018e-08
Rx480 x480 0 1
Fxc480_479 x480 0 Vx479 -1172.08639744215
Cx480 x480 xm480 6.6456706498173e-14
Vx480 xm480 0 0
Gx480_1 x480 0 u1 0 3.37385051730226e-05
Rx481 x481 0 1
Fxc481_482 x481 0 Vx482 33.9357310812671
Cx481 x481 xm481 1.92779692469307e-13
Vx481 xm481 0 0
Gx481_1 x481 0 u1 0 -8.83869563481327e-08
Rx482 x482 0 1
Fxc482_481 x482 0 Vx481 -1235.73548395772
Cx482 x482 xm482 1.92779692469307e-13
Vx482 xm482 0 0
Gx482_1 x482 0 u1 0 0.00010922289827841
Rx483 x483 0 1
Fxc483_484 x483 0 Vx484 261.34138678253
Cx483 x483 xm483 1.15282449142532e-12
Vx483 xm483 0 0
Gx483_1 x483 0 u1 0 -9.8275060838972e-05
Rx484 x484 0 1
Fxc484_483 x484 0 Vx483 -4.99147261695213
Cx484 x484 xm484 1.15282449142532e-12
Vx484 xm484 0 0
Gx484_1 x484 0 u1 0 0.000490537275107034
Rx485 x485 0 1
Fxc485_486 x485 0 Vx486 9688.80562447404
Cx485 x485 xm485 2.87628016359056e-14
Vx485 xm485 0 0
Gx485_1 x485 0 u1 0 -3.94315662075411e-09
Rx486 x486 0 1
Fxc486_485 x486 0 Vx485 -195.064678811955
Cx486 x486 xm486 2.87628016359056e-14
Vx486 xm486 0 0
Gx486_1 x486 0 u1 0 7.69170579732633e-07
Rx487 x487 0 1
Fxc487_488 x487 0 Vx488 22.9370756708558
Cx487 x487 xm487 1.78666875824597e-13
Vx487 xm487 0 0
Gx487_1 x487 0 u1 0 -5.73359517242577e-08
Rx488 x488 0 1
Fxc488_487 x488 0 Vx487 -2184.16581406027
Cx488 x488 xm488 1.78666875824597e-13
Vx488 xm488 0 0
Gx488_1 x488 0 u1 0 0.000125231225672734
Rx489 x489 0 1
Fxc489_490 x489 0 Vx490 1333.40746689041
Cx489 x489 xm489 1.04155247034917e-13
Vx489 xm489 0 0
Gx489_1 x489 0 u1 0 -1.34649883907356e-07
Rx490 x490 0 1
Fxc490_489 x490 0 Vx489 -109.715007510101
Cx490 x490 xm490 1.04155247034917e-13
Vx490 xm490 0 0
Gx490_1 x490 0 u1 0 1.47731130241297e-05
Rx491 x491 0 1
Fxc491_492 x491 0 Vx492 926.132810904575
Cx491 x491 xm491 1.06235443062179e-14
Vx491 xm491 0 0
Gx491_1 x491 0 u1 0 -3.71468040427725e-10
Rx492 x492 0 1
Fxc492_491 x492 0 Vx491 -15597.5586059317
Cx492 x492 xm492 1.06235443062179e-14
Vx492 xm492 0 0
Gx492_1 x492 0 u1 0 5.79399453080205e-06
Rx493 x493 0 1
Fxc493_494 x493 0 Vx494 353.970852756558
Cx493 x493 xm493 5.41238890095385e-14
Vx493 xm493 0 0
Gx493_1 x493 0 u1 0 -7.06659962780316e-09
Rx494 x494 0 1
Fxc494_493 x494 0 Vx493 -1599.44081251103
Cx494 x494 xm494 5.41238890095385e-14
Vx494 xm494 0 0
Gx494_1 x494 0 u1 0 1.13026078503837e-05
Rx495 x495 0 1
Fxc495_496 x495 0 Vx496 2390.13634534209
Cx495 x495 xm495 3.3864832840636e-14
Vx495 xm495 0 0
Gx495_1 x495 0 u1 0 -8.6055070507376e-09
Rx496 x496 0 1
Fxc496_495 x496 0 Vx495 -611.532670584081
Cx496 x496 xm496 3.3864832840636e-14
Vx496 xm496 0 0
Gx496_1 x496 0 u1 0 5.2625487084677e-06
Rx497 x497 0 1
Fxc497_498 x497 0 Vx498 35.945069362476
Cx497 x497 xm497 4.1684778621004e-13
Vx497 xm497 0 0
Gx497_1 x497 0 u1 0 -2.14315186580318e-06
Rx498 x498 0 1
Fxc498_497 x498 0 Vx497 -282.624295333059
Cx498 x498 xm498 4.1684778621004e-13
Vx498 xm498 0 0
Gx498_1 x498 0 u1 0 0.000605706785864354
Rx499 x499 0 1
Fxc499_500 x499 0 Vx500 996.665715892896
Cx499 x499 xm499 1.43290144219323e-14
Vx499 xm499 0 0
Gx499_1 x499 0 u1 0 -9.13742982859077e-10
Rx500 x500 0 1
Fxc500_499 x500 0 Vx499 -8387.30918589729
Cx500 x500 xm500 1.43290144219323e-14
Vx500 xm500 0 0
Gx500_1 x500 0 u1 0 7.66384491368313e-06
Rx501 x501 0 1
Fxc501_502 x501 0 Vx502 918.277931646278
Cx501 x501 xm501 1.59153780242877e-14
Vx501 xm501 0 0
Gx501_1 x501 0 u1 0 -1.26635722230678e-09
Rx502 x502 0 1
Fxc502_501 x502 0 Vx501 -7843.21116664781
Cx502 x502 xm502 1.59153780242877e-14
Vx502 xm502 0 0
Gx502_1 x502 0 u1 0 9.93230710696161e-06
Rx503 x503 0 1
Fxc503_504 x503 0 Vx504 1314.17217114326
Cx503 x503 xm503 1.1293667793922e-13
Vx503 xm503 0 0
Gx503_1 x503 0 u1 0 -6.3622907491661e-08
Rx504 x504 0 1
Fxc504_503 x504 0 Vx503 -107.870021691714
Cx504 x504 xm504 1.1293667793922e-13
Vx504 xm504 0 0
Gx504_1 x504 0 u1 0 6.86300441121535e-06
Rx505 x505 0 1
Fxc505_506 x505 0 Vx506 441.219514187201
Cx505 x505 xm505 1.00794993851598e-13
Vx505 xm505 0 0
Gx505_1 x505 0 u1 0 -7.88094719322437e-08
Rx506 x506 0 1
Fxc506_505 x506 0 Vx505 -397.404591516267
Cx506 x506 xm506 1.00794993851598e-13
Vx506 xm506 0 0
Gx506_1 x506 0 u1 0 3.1319246000846e-05
Rx507 x507 0 1
Fxc507_508 x507 0 Vx508 453.700505163878
Cx507 x507 xm507 3.93436377555167e-14
Vx507 xm507 0 0
Gx507_1 x507 0 u1 0 -5.50907702795513e-09
Rx508 x508 0 1
Fxc508_507 x508 0 Vx507 -2503.33256649344
Cx508 x508 xm508 3.93436377555167e-14
Vx508 xm508 0 0
Gx508_1 x508 0 u1 0 1.3791051935401e-05
Rx509 x509 0 1
Fxc509_510 x509 0 Vx510 1565.23641201402
Cx509 x509 xm509 4.27323643580748e-14
Vx509 xm509 0 0
Gx509_1 x509 0 u1 0 -3.20532174022322e-09
Rx510 x510 0 1
Fxc510_509 x510 0 Vx509 -653.806833195912
Cx510 x510 xm510 4.27323643580748e-14
Vx510 xm510 0 0
Gx510_1 x510 0 u1 0 2.09566125634935e-06
Rx511 x511 0 1
Cx511 x511 0 1.40144076963712e-10
Gx511_1 x511 0 u1 0 -9.91549848804308
Rx512 x512 0 1
Fxc512_513 x512 0 Vx513 40.9099257192964
Cx512 x512 xm512 1.39431711841145e-12
Vx512 xm512 0 0
Gx512_1 x512 0 u1 0 -0.000159753606995055
Rx513 x513 0 1
Fxc513_512 x513 0 Vx512 -27.1610623814526
Cx513 x513 xm513 1.39431711841145e-12
Vx513 xm513 0 0
Gx513_1 x513 0 u1 0 0.00433907768525475
Rx514 x514 0 1
Fxc514_515 x514 0 Vx515 1271.99120570634
Cx514 x514 xm514 4.46055376469595e-14
Vx514 xm514 0 0
Gx514_1 x514 0 u1 0 -7.90118001768697e-09
Rx515 x515 0 1
Fxc515_514 x515 0 Vx514 -813.486312276597
Cx515 x515 xm515 4.46055376469595e-14
Vx515 xm515 0 0
Gx515_1 x515 0 u1 0 6.42750179522171e-06
Rx516 x516 0 1
Fxc516_517 x516 0 Vx517 386.18834089681
Cx516 x516 xm516 1.38311295911203e-13
Vx516 xm516 0 0
Gx516_1 x516 0 u1 0 -4.07163779962862e-07
Rx517 x517 0 1
Fxc517_516 x517 0 Vx516 -269.303864140825
Cx517 x517 xm517 1.38311295911203e-13
Vx517 xm517 0 0
Gx517_1 x517 0 u1 0 0.000109650779282183
Rx518 x518 0 1
Fxc518_519 x518 0 Vx519 76.2968719363534
Cx518 x518 xm518 2.19578957008743e-13
Vx518 xm518 0 0
Gx518_1 x518 0 u1 0 -5.94382313711905e-07
Rx519 x519 0 1
Fxc519_518 x519 0 Vx518 -541.968774581695
Cx519 x519 xm519 2.19578957008743e-13
Vx519 xm519 0 0
Gx519_1 x519 0 u1 0 0.000322136654195474
Rx520 x520 0 1
Fxc520_521 x520 0 Vx521 842.159723820827
Cx520 x520 xm520 4.73505553997717e-14
Vx520 xm520 0 0
Gx520_1 x520 0 u1 0 -9.34487758818243e-09
Rx521 x521 0 1
Fxc521_520 x521 0 Vx520 -1010.88481543308
Cx521 x521 xm521 4.73505553997717e-14
Vx521 xm521 0 0
Gx521_1 x521 0 u1 0 9.44659485597452e-06
Rx522 x522 0 1
Fxc522_523 x522 0 Vx523 115.364127646596
Cx522 x522 xm522 1.22056182242707e-13
Vx522 xm522 0 0
Gx522_1 x522 0 u1 0 -4.63136413714817e-08
Rx523 x523 0 1
Fxc523_522 x523 0 Vx522 -1124.95887344488
Cx523 x523 xm523 1.22056182242707e-13
Vx523 xm523 0 0
Gx523_1 x523 0 u1 0 5.21009418223923e-05
Rx524 x524 0 1
Fxc524_525 x524 0 Vx525 657.85532305545
Cx524 x524 xm524 4.2540439057887e-14
Vx524 xm524 0 0
Gx524_1 x524 0 u1 0 -9.38487669122894e-09
Rx525 x525 0 1
Fxc525_524 x525 0 Vx524 -1646.38526251394
Cx525 x525 xm525 4.2540439057887e-14
Vx525 xm525 0 0
Gx525_1 x525 0 u1 0 1.54511226749499e-05
Rx526 x526 0 1
Fxc526_527 x526 0 Vx527 0.605110726296806
Cx526 x526 xm526 8.16769439323924e-11
Vx526 xm526 0 0
Gx526_1 x526 0 u1 0 -4.69783978368822
Rx527 x527 0 1
Fxc527_526 x527 0 Vx526 -1.12450076992043
Cx527 x527 xm527 8.16769439323924e-11
Vx527 xm527 0 0
Gx527_1 x527 0 u1 0 5.28272445372025
Rx528 x528 0 1
Fxc528_529 x528 0 Vx529 2.21091652567028
Cx528 x528 xm528 3.055355601781e-12
Vx528 xm528 0 0
Gx528_1 x528 0 u1 0 -0.000185389851087876
Rx529 x529 0 1
Fxc529_528 x529 0 Vx528 -119.071455429122
Cx529 x529 xm529 3.055355601781e-12
Vx529 xm529 0 0
Gx529_1 x529 0 u1 0 0.0220746393908216
Rx530 x530 0 1
Fxc530_531 x530 0 Vx531 95.2035374767698
Cx530 x530 xm530 2.22336076590458e-13
Vx530 xm530 0 0
Gx530_1 x530 0 u1 0 -2.3985141742488e-07
Rx531 x531 0 1
Fxc531_530 x531 0 Vx530 -524.093472474892
Cx531 x531 xm531 2.22336076590458e-13
Vx531 xm531 0 0
Gx531_1 x531 0 u1 0 0.00012570456223623
Rx532 x532 0 1
Fxc532_533 x532 0 Vx533 52.6156141590728
Cx532 x532 xm532 7.0682437690172e-13
Vx532 xm532 0 0
Gx532_1 x532 0 u1 0 -1.55913839594535e-05
Rx533 x533 0 1
Fxc533_532 x533 0 Vx532 -84.9724515057839
Cx533 x533 xm533 7.0682437690172e-13
Vx533 xm533 0 0
Gx533_1 x533 0 u1 0 0.00132483811740272
Rx534 x534 0 1
Fxc534_535 x534 0 Vx535 1108.20901796368
Cx534 x534 xm534 5.1045195384584e-14
Vx534 xm534 0 0
Gx534_1 x534 0 u1 0 -9.44918798334939e-09
Rx535 x535 0 1
Fxc535_534 x535 0 Vx534 -724.595992548357
Cx535 x535 xm535 5.1045195384584e-14
Vx535 xm535 0 0
Gx535_1 x535 0 u1 0 6.84684374557106e-06
Rx536 x536 0 1
Fxc536_537 x536 0 Vx537 1942.43973474849
Cx536 x536 xm536 2.41223264060163e-13
Vx536 xm536 0 0
Gx536_1 x536 0 u1 0 -5.7707596304258e-07
Rx537 x537 0 1
Fxc537_536 x537 0 Vx536 -18.9908482522893
Cx537 x537 xm537 2.41223264060163e-13
Vx537 xm537 0 0
Gx537_1 x537 0 u1 0 1.09591620441853e-05
Rx538 x538 0 1
Fxc538_539 x538 0 Vx539 1308.30023135288
Cx538 x538 xm538 9.93476076097149e-14
Vx538 xm538 0 0
Gx538_1 x538 0 u1 0 -5.71496833314397e-08
Rx539 x539 0 1
Fxc539_538 x539 0 Vx538 -168.785335337332
Cx539 x539 xm539 9.93476076097149e-14
Vx539 xm539 0 0
Gx539_1 x539 0 u1 0 9.64602846551938e-06
Rx540 x540 0 1
Fxc540_541 x540 0 Vx541 289.041515254048
Cx540 x540 xm540 1.96255535649835e-14
Vx540 xm540 0 0
Gx540_1 x540 0 u1 0 -8.08009149132606e-10
Rx541 x541 0 1
Fxc541_540 x541 0 Vx540 -20108.7876320356
Cx541 x541 xm541 1.96255535649835e-14
Vx541 xm541 0 0
Gx541_1 x541 0 u1 0 1.62480843846493e-05
Rx542 x542 0 1
Fxc542_543 x542 0 Vx543 268.465853463582
Cx542 x542 xm542 2.15369618623669e-13
Vx542 xm542 0 0
Gx542_1 x542 0 u1 0 -3.25800201565287e-07
Rx543 x543 0 1
Fxc543_542 x543 0 Vx542 -184.48774922061
Cx543 x543 xm543 2.15369618623669e-13
Vx543 xm543 0 0
Gx543_1 x543 0 u1 0 6.0106145882401e-05
Rx544 x544 0 1
Fxc544_545 x544 0 Vx545 1138.40970836513
Cx544 x544 xm544 1.21891798583539e-14
Vx544 xm544 0 0
Gx544_1 x544 0 u1 0 -1.86273421242884e-10
Rx545 x545 0 1
Fxc545_544 x545 0 Vx544 -12532.3923557284
Cx545 x545 xm545 1.21891798583539e-14
Vx545 xm545 0 0
Gx545_1 x545 0 u1 0 2.33445160045969e-06
Rx546 x546 0 1
Fxc546_547 x546 0 Vx547 5244.27905038958
Cx546 x546 xm546 2.69942236556942e-14
Vx546 xm546 0 0
Gx546_1 x546 0 u1 0 -5.97906372382909e-09
Rx547 x547 0 1
Fxc547_546 x547 0 Vx546 -630.461550836563
Cx547 x547 xm547 2.69942236556942e-14
Vx547 xm547 0 0
Gx547_1 x547 0 u1 0 3.76956978787593e-06
Rx548 x548 0 1
Fxc548_549 x548 0 Vx549 23.8525173809244
Cx548 x548 xm548 7.7544284673081e-14
Vx548 xm548 0 0
Gx548_1 x548 0 u1 0 -1.05252836908603e-09
Rx549 x549 0 1
Fxc549_548 x549 0 Vx548 -16290.2204910886
Cx549 x549 xm549 7.7544284673081e-14
Vx549 xm549 0 0
Gx549_1 x549 0 u1 0 1.71459192055373e-05
Rx550 x550 0 1
Fxc550_551 x550 0 Vx551 1022.86453608461
Cx550 x550 xm550 1.03543939234814e-13
Vx550 xm550 0 0
Gx550_1 x550 0 u1 0 -5.69665671548081e-08
Rx551 x551 0 1
Fxc551_550 x551 0 Vx550 -216.837694283884
Cx551 x551 xm551 1.03543939234814e-13
Vx551 xm551 0 0
Gx551_1 x551 0 u1 0 1.23524990731166e-05
Rx552 x552 0 1
Fxc552_553 x552 0 Vx553 781.237041345032
Cx552 x552 xm552 9.1674395278034e-14
Vx552 xm552 0 0
Gx552_1 x552 0 u1 0 -5.68790784729225e-08
Rx553 x553 0 1
Fxc553_552 x553 0 Vx552 -378.142571801365
Cx553 x553 xm553 9.1674395278034e-14
Vx553 xm553 0 0
Gx553_1 x553 0 u1 0 2.15084010154425e-05
Rx554 x554 0 1
Fxc554_555 x554 0 Vx555 153.311464854679
Cx554 x554 xm554 1.90368710342961e-13
Vx554 xm554 0 0
Gx554_1 x554 0 u1 0 -1.06843518202555e-07
Rx555 x555 0 1
Fxc555_554 x555 0 Vx554 -461.4522145074
Cx555 x555 xm555 1.90368710342961e-13
Vx555 xm555 0 0
Gx555_1 x555 0 u1 0 4.93031780803309e-05
Rx556 x556 0 1
Fxc556_557 x556 0 Vx557 13802.952547307
Cx556 x556 xm556 3.43839976006569e-14
Vx556 xm556 0 0
Gx556_1 x556 0 u1 0 -3.21278576409548e-09
Rx557 x557 0 1
Fxc557_556 x557 0 Vx556 -158.289370739167
Cx557 x557 xm557 3.43839976006569e-14
Vx557 xm557 0 0
Gx557_1 x557 0 u1 0 5.08549836918429e-07
Rx558 x558 0 1
Fxc558_559 x558 0 Vx559 2449.36498759504
Cx558 x558 xm558 1.10377999804161e-13
Vx558 xm558 0 0
Gx558_1 x558 0 u1 0 -2.63022165275067e-08
Rx559 x559 0 1
Fxc559_558 x559 0 Vx558 -87.9776222078131
Cx559 x559 xm559 1.10377999804161e-13
Vx559 xm559 0 0
Gx559_1 x559 0 u1 0 2.31400646888508e-06
Rx560 x560 0 1
Fxc560_561 x560 0 Vx561 13419.594844209
Cx560 x560 xm560 5.39843163452879e-14
Vx560 xm560 0 0
Gx560_1 x560 0 u1 0 -1.14009821937492e-08
Rx561 x561 0 1
Fxc561_560 x561 0 Vx560 -68.936724154623
Cx561 x561 xm561 5.39843163452879e-14
Vx561 xm561 0 0
Gx561_1 x561 0 u1 0 7.85946364582258e-07
Rx562 x562 0 1
Fxc562_563 x562 0 Vx563 929.96862403055
Cx562 x562 xm562 1.66115615183985e-13
Vx562 xm562 0 0
Gx562_1 x562 0 u1 0 -1.62146499736644e-07
Rx563 x563 0 1
Fxc563_562 x563 0 Vx562 -106.633817486013
Cx563 x563 xm563 1.66115615183985e-13
Vx563 xm563 0 0
Gx563_1 x563 0 u1 0 1.72903002589133e-05
Rx564 x564 0 1
Fxc564_565 x564 0 Vx565 23123.4177217671
Cx564 x564 xm564 1.72753550245707e-13
Vx564 xm564 0 0
Gx564_1 x564 0 u1 0 -7.31080462978585e-07
Rx565 x565 0 1
Fxc565_564 x565 0 Vx564 -4.0530113543923
Cx565 x565 xm565 1.72753550245707e-13
Vx565 xm565 0 0
Gx565_1 x565 0 u1 0 2.96307741742658e-06
Rx566 x566 0 1
Fxc566_567 x566 0 Vx567 3086.48100565301
Cx566 x566 xm566 7.89077374985022e-14
Vx566 xm566 0 0
Gx566_1 x566 0 u1 0 -1.20816551927519e-07
Rx567 x567 0 1
Fxc567_566 x567 0 Vx566 -145.44136304278
Cx567 x567 xm567 7.89077374985022e-14
Vx567 xm567 0 0
Gx567_1 x567 0 u1 0 1.75717239904673e-05
Rx568 x568 0 1
Fxc568_569 x568 0 Vx569 78.8366728598425
Cx568 x568 xm568 4.41676639181862e-13
Vx568 xm568 0 0
Gx568_1 x568 0 u1 0 -3.25901533117844e-06
Rx569 x569 0 1
Fxc569_568 x569 0 Vx568 -187.227487667191
Cx569 x569 xm569 4.41676639181862e-13
Vx569 xm569 0 0
Gx569_1 x569 0 u1 0 0.000610177252725399
Rx570 x570 0 1
Fxc570_571 x570 0 Vx571 90.843312542467
Cx570 x570 xm570 7.69508360165092e-13
Vx570 xm570 0 0
Gx570_1 x570 0 u1 0 -8.66949332050594e-05
Rx571 x571 0 1
Fxc571_570 x571 0 Vx570 -55.5692884423165
Cx571 x571 xm571 7.69508360165092e-13
Vx571 xm571 0 0
Gx571_1 x571 0 u1 0 0.00481757574975931
Rx572 x572 0 1
Fxc572_573 x572 0 Vx573 2907.73543531577
Cx572 x572 xm572 6.84174064919173e-13
Vx572 xm572 0 0
Gx572_1 x572 0 u1 0 -0.000117312262866649
Rx573 x573 0 1
Fxc573_572 x573 0 Vx572 -2.17266166295278
Cx573 x573 xm573 6.84174064919173e-13
Vx573 xm573 0 0
Gx573_1 x573 0 u1 0 0.000254879856124608
Rx574 x574 0 1
Fxc574_575 x574 0 Vx575 5830.55830943377
Cx574 x574 xm574 3.41606667996328e-13
Vx574 xm574 0 0
Gx574_1 x574 0 u1 0 -5.97471694796694e-06
Rx575 x575 0 1
Fxc575_574 x575 0 Vx574 -4.33839407522684
Cx575 x575 xm575 3.41606667996328e-13
Vx575 xm575 0 0
Gx575_1 x575 0 u1 0 2.59206766082171e-05
Rx576 x576 0 1
Fxc576_577 x576 0 Vx577 20.1556839267652
Cx576 x576 xm576 1.07548830475537e-12
Vx576 xm576 0 0
Gx576_1 x576 0 u1 0 -1.50845268902827e-05
Rx577 x577 0 1
Fxc577_576 x577 0 Vx576 -135.904079368811
Cx577 x577 xm577 1.07548830475537e-12
Vx577 xm577 0 0
Gx577_1 x577 0 u1 0 0.00205004873973794
Rx578 x578 0 1
Fxc578_579 x578 0 Vx579 160.732494484157
Cx578 x578 xm578 1.99049200010659e-13
Vx578 xm578 0 0
Gx578_1 x578 0 u1 0 -1.00004422141991e-07
Rx579 x579 0 1
Fxc579_578 x579 0 Vx578 -499.319998397926
Cx579 x579 xm579 1.99049200010659e-13
Vx579 xm579 0 0
Gx579_1 x579 0 u1 0 4.99342079037243e-05
Rx580 x580 0 1
Fxc580_581 x580 0 Vx581 150.576720409034
Cx580 x580 xm580 1.88237358199619e-13
Vx580 xm580 0 0
Gx580_1 x580 0 u1 0 -8.1470253881492e-08
Rx581 x581 0 1
Fxc581_580 x581 0 Vx580 -577.741724916063
Cx581 x581 xm581 1.88237358199619e-13
Vx581 xm581 0 0
Gx581_1 x581 0 u1 0 4.70687650068427e-05
Rx582 x582 0 1
Fxc582_583 x582 0 Vx583 22958.4508175614
Cx582 x582 xm582 1.57459489839352e-14
Vx582 xm582 0 0
Gx582_1 x582 0 u1 0 -6.65923190185912e-10
Rx583 x583 0 1
Fxc583_582 x583 0 Vx582 -531.225813529373
Cx583 x583 xm583 1.57459489839352e-14
Vx583 xm583 0 0
Gx583_1 x583 0 u1 0 3.53755588454587e-07
Rx584 x584 0 1
Fxc584_585 x584 0 Vx585 2683.91607243587
Cx584 x584 xm584 2.49001986220754e-14
Vx584 xm584 0 0
Gx584_1 x584 0 u1 0 -1.36801420560313e-09
Rx585 x585 0 1
Fxc585_584 x585 0 Vx584 -2039.16542494762
Cx585 x585 xm585 2.49001986220754e-14
Vx585 xm585 0 0
Gx585_1 x585 0 u1 0 2.78960726890308e-06
Rx586 x586 0 1
Fxc586_587 x586 0 Vx587 49.6224004425067
Cx586 x586 xm586 1.20010327111104e-13
Vx586 xm586 0 0
Gx586_1 x586 0 u1 0 -4.60410846045463e-09
Rx587 x587 0 1
Fxc587_586 x587 0 Vx586 -4637.77693820943
Cx587 x587 xm587 1.20010327111104e-13
Vx587 xm587 0 0
Gx587_1 x587 0 u1 0 2.13528280389114e-05
Rx588 x588 0 1
Fxc588_589 x588 0 Vx589 113.680054486503
Cx588 x588 xm588 9.19589919698257e-13
Vx588 xm588 0 0
Gx588_1 x588 0 u1 0 -3.67918786745731e-05
Rx589 x589 0 1
Fxc589_588 x589 0 Vx588 -37.0988060597012
Cx589 x589 xm589 9.19589919698257e-13
Vx589 xm589 0 0
Gx589_1 x589 0 u1 0 0.00136493477152005
Rx590 x590 0 1
Fxc590_591 x590 0 Vx591 92.5261479237949
Cx590 x590 xm590 1.35062615998325e-12
Vx590 xm590 0 0
Gx590_1 x590 0 u1 0 -0.000130795948893988
Rx591 x591 0 1
Fxc591_590 x591 0 Vx590 -21.1941138098059
Cx591 x591 xm591 1.35062615998325e-12
Vx591 xm591 0 0
Gx591_1 x591 0 u1 0 0.00277210422672074
Rx592 x592 0 1
Fxc592_593 x592 0 Vx593 18792.6439027955
Cx592 x592 xm592 5.61403593569498e-16
Vx592 xm592 0 0
Gx592_1 x592 0 u1 0 -1.23966122217621e-11
Rx593 x593 0 1
Fxc593_592 x593 0 Vx592 -590684.859353706
Cx593 x593 xm593 5.61403593569498e-16
Vx593 xm593 0 0
Gx593_1 x593 0 u1 0 7.32249114667396e-06
Rx594 x594 0 1
Fxc594_595 x594 0 Vx595 264.99743569509
Cx594 x594 xm594 1.34555540326277e-13
Vx594 xm594 0 0
Gx594_1 x594 0 u1 0 -4.23658539188337e-08
Rx595 x595 0 1
Fxc595_594 x595 0 Vx594 -749.798059430211
Cx595 x595 xm595 1.34555540326277e-13
Vx595 xm595 0 0
Gx595_1 x595 0 u1 0 3.17658350544453e-05
Rx596 x596 0 1
Fxc596_597 x596 0 Vx597 690.978884695212
Cx596 x596 xm596 4.98865404960471e-13
Vx596 xm596 0 0
Gx596_1 x596 0 u1 0 -1.66025322113517e-06
Rx597 x597 0 1
Fxc597_596 x597 0 Vx596 -25.4811031218623
Cx597 x597 xm597 4.98865404960471e-13
Vx597 xm597 0 0
Gx597_1 x597 0 u1 0 4.23050835361492e-05
Rx598 x598 0 1
Fxc598_599 x598 0 Vx599 75.9454614588599
Cx598 x598 xm598 1.15714797739341e-12
Vx598 xm598 0 0
Gx598_1 x598 0 u1 0 -2.07458779796158e-05
Rx599 x599 0 1
Fxc599_598 x599 0 Vx598 -38.2863285868415
Cx599 x599 xm599 1.15714797739341e-12
Vx599 xm599 0 0
Gx599_1 x599 0 u1 0 0.000794283501150088
Rx600 x600 0 1
Fxc600_601 x600 0 Vx601 82.2567761245647
Cx600 x600 xm600 5.42048534221595e-13
Vx600 xm600 0 0
Gx600_1 x600 0 u1 0 -1.91865879274409e-06
Rx601 x601 0 1
Fxc601_600 x601 0 Vx600 -169.803176527306
Cx601 x601 xm601 5.42048534221595e-13
Vx601 xm601 0 0
Gx601_1 x601 0 u1 0 0.000325794357679993
Rx602 x602 0 1
Fxc602_603 x602 0 Vx603 917.827176623362
Cx602 x602 xm602 9.340099268043e-14
Vx602 xm602 0 0
Gx602_1 x602 0 u1 0 -1.4095703771799e-08
Rx603 x603 0 1
Fxc603_602 x603 0 Vx602 -474.731753891079
Cx603 x603 xm603 9.340099268043e-14
Vx603 xm603 0 0
Gx603_1 x603 0 u1 0 6.69167817391524e-06
Rx604 x604 0 1
Fxc604_605 x604 0 Vx605 358.739707000422
Cx604 x604 xm604 2.02797650128333e-13
Vx604 xm604 0 0
Gx604_1 x604 0 u1 0 -1.00673054246152e-07
Rx605 x605 0 1
Fxc605_604 x605 0 Vx604 -285.960066242383
Cx605 x605 xm605 2.02797650128333e-13
Vx605 xm605 0 0
Gx605_1 x605 0 u1 0 2.87884732610527e-05
Rx606 x606 0 1
Fxc606_607 x606 0 Vx607 90.1170888923772
Cx606 x606 xm606 7.01742537232251e-13
Vx606 xm606 0 0
Gx606_1 x606 0 u1 0 -6.15344149099034e-06
Rx607 x607 0 1
Fxc607_606 x607 0 Vx606 -93.7539039129234
Cx607 x607 xm607 7.01742537232251e-13
Vx607 xm607 0 0
Gx607_1 x607 0 u1 0 0.000576909162280105
Rx608 x608 0 1
Fxc608_609 x608 0 Vx609 613.253330633679
Cx608 x608 xm608 6.4028082506253e-14
Vx608 xm608 0 0
Gx608_1 x608 0 u1 0 -7.83594578363736e-09
Rx609 x609 0 1
Fxc609_608 x609 0 Vx608 -1479.08238714529
Cx609 x609 xm609 6.4028082506253e-14
Vx609 xm609 0 0
Gx609_1 x609 0 u1 0 1.15900093952034e-05
Rx610 x610 0 1
Fxc610_611 x610 0 Vx611 6557.81169373482
Cx610 x610 xm610 3.68280434719191e-14
Vx610 xm610 0 0
Gx610_1 x610 0 u1 0 -4.23599676313272e-09
Rx611 x611 0 1
Fxc611_610 x611 0 Vx610 -446.872773418864
Cx611 x611 xm611 3.68280434719191e-14
Vx611 xm611 0 0
Gx611_1 x611 0 u1 0 1.89295162173445e-06
Rx612 x612 0 1
Fxc612_613 x612 0 Vx613 319.312683895813
Cx612 x612 xm612 2.43463431944243e-13
Vx612 xm612 0 0
Gx612_1 x612 0 u1 0 -1.57458933118466e-07
Rx613 x613 0 1
Fxc613_612 x613 0 Vx612 -202.786593577218
Cx613 x613 xm613 2.43463431944243e-13
Vx613 xm613 0 0
Gx613_1 x613 0 u1 0 3.19305606753967e-05
Rx614 x614 0 1
Fxc614_615 x614 0 Vx615 1489.29144013567
Cx614 x614 xm614 1.88338702913179e-13
Vx614 xm614 0 0
Gx614_1 x614 0 u1 0 -1.03956884002395e-07
Rx615 x615 0 1
Fxc615_614 x615 0 Vx614 -82.9218259369898
Cx615 x615 xm615 1.88338702913179e-13
Vx615 xm615 0 0
Gx615_1 x615 0 u1 0 8.62029464019842e-06
Rx616 x616 0 1
Fxc616_617 x616 0 Vx617 16191.1108915013
Cx616 x616 xm616 4.99523803066435e-15
Vx616 xm616 0 0
Gx616_1 x616 0 u1 0 -7.41077976107855e-10
Rx617 x617 0 1
Fxc617_616 x617 0 Vx616 -11188.052581356
Cx617 x617 xm617 4.99523803066435e-15
Vx617 xm617 0 0
Gx617_1 x617 0 u1 0 8.29121936357956e-06
Rx618 x618 0 1
Fxc618_619 x618 0 Vx619 0.820660349771105
Cx618 x618 xm618 7.43266824125504e-12
Vx618 xm618 0 0
Gx618_1 x618 0 u1 0 -0.000648728921442811
Rx619 x619 0 1
Fxc619_618 x619 0 Vx618 -130.604943847461
Cx619 x619 xm619 7.43266824125504e-12
Vx619 xm619 0 0
Gx619_1 x619 0 u1 0 0.0847272043572624
Rx620 x620 0 1
Fxc620_621 x620 0 Vx621 35.6681472841325
Cx620 x620 xm620 1.3706119903344e-12
Vx620 xm620 0 0
Gx620_1 x620 0 u1 0 -8.83398825978201e-06
Rx621 x621 0 1
Fxc621_620 x621 0 Vx620 -72.2604353179937
Cx621 x621 xm621 1.3706119903344e-12
Vx621 xm621 0 0
Gx621_1 x621 0 u1 0 0.000638347837245893
Rx622 x622 0 1
Fxc622_623 x622 0 Vx623 4519.69639650926
Cx622 x622 xm622 1.32600732830319e-13
Vx622 xm622 0 0
Gx622_1 x622 0 u1 0 -3.05308186797716e-08
Rx623 x623 0 1
Fxc623_622 x623 0 Vx622 -59.6341007177601
Cx623 x623 xm623 1.32600732830319e-13
Vx623 xm623 0 0
Gx623_1 x623 0 u1 0 1.82067791614517e-06
Rx624 x624 0 1
Fxc624_625 x624 0 Vx625 1313.10638550444
Cx624 x624 xm624 6.7800124285245e-14
Vx624 xm624 0 0
Gx624_1 x624 0 u1 0 -1.37489855025595e-08
Rx625 x625 0 1
Fxc625_624 x625 0 Vx624 -809.411391209405
Cx625 x625 xm625 6.7800124285245e-14
Vx625 xm625 0 0
Gx625_1 x625 0 u1 0 1.11285854833446e-05
Rx626 x626 0 1
Fxc626_627 x626 0 Vx627 218.814403501971
Cx626 x626 xm626 1.115641621969e-13
Vx626 xm626 0 0
Gx626_1 x626 0 u1 0 -1.27488894192533e-08
Rx627 x627 0 1
Fxc627_626 x627 0 Vx626 -1833.28842657534
Cx627 x627 xm627 1.115641621969e-13
Vx627 xm627 0 0
Gx627_1 x627 0 u1 0 2.33723914240058e-05
Rx628 x628 0 1
Fxc628_629 x628 0 Vx629 66.1480927412148
Cx628 x628 xm628 2.72702074238325e-13
Vx628 xm628 0 0
Gx628_1 x628 0 u1 0 -3.69778853644285e-08
Rx629 x629 0 1
Fxc629_628 x629 0 Vx628 -1062.7570648512
Cx629 x629 xm629 2.72702074238325e-13
Vx629 xm629 0 0
Gx629_1 x629 0 u1 0 3.92985089143042e-05
Rx630 x630 0 1
Fxc630_631 x630 0 Vx631 39.5010738646823
Cx630 x630 xm630 1.01079656034734e-12
Vx630 xm630 0 0
Gx630_1 x630 0 u1 0 -4.9715514735905e-06
Rx631 x631 0 1
Fxc631_630 x631 0 Vx630 -134.429386049206
Cx631 x631 xm631 1.01079656034734e-12
Vx631 xm631 0 0
Gx631_1 x631 0 u1 0 0.000668322612306796
Rx632 x632 0 1
Fxc632_633 x632 0 Vx633 1344.06085477589
Cx632 x632 xm632 8.24832104280923e-14
Vx632 xm632 0 0
Gx632_1 x632 0 u1 0 -1.86132702602691e-08
Rx633 x633 0 1
Fxc633_632 x633 0 Vx632 -582.660599826319
Cx633 x633 xm633 8.24832104280923e-14
Vx633 xm633 0 0
Gx633_1 x633 0 u1 0 1.08452192145778e-05
Rx634 x634 0 1
Fxc634_635 x634 0 Vx635 607.733912981475
Cx634 x634 xm634 2.39433153810415e-13
Vx634 xm634 0 0
Gx634_1 x634 0 u1 0 -1.36276240736005e-07
Rx635 x635 0 1
Fxc635_634 x635 0 Vx634 -157.939337993207
Cx635 x635 xm635 2.39433153810415e-13
Vx635 xm635 0 0
Gx635_1 x635 0 u1 0 2.15233792460475e-05
Rx636 x636 0 1
Fxc636_637 x636 0 Vx637 23.2940179636851
Cx636 x636 xm636 2.46268600071512e-12
Vx636 xm636 0 0
Gx636_1 x636 0 u1 0 -0.000411254870970819
Rx637 x637 0 1
Fxc637_636 x637 0 Vx636 -44.2825934935633
Cx637 x637 xm637 2.46268600071512e-12
Vx637 xm637 0 0
Gx637_1 x637 0 u1 0 0.0182114322734486
Rx638 x638 0 1
Fxc638_639 x638 0 Vx639 14.0841777848976
Cx638 x638 xm638 3.96234308451515e-12
Vx638 xm638 0 0
Gx638_1 x638 0 u1 0 -0.00016473305947621
Rx639 x639 0 1
Fxc639_638 x639 0 Vx638 -36.1159740107871
Cx639 x639 xm639 3.96234308451514e-12
Vx639 xm639 0 0
Gx639_1 x639 0 u1 0 0.00594949489476025
Rx640 x640 0 1
Fxc640_641 x640 0 Vx641 1086.43095441727
Cx640 x640 xm640 8.60345839298812e-13
Vx640 xm640 0 0
Gx640_1 x640 0 u1 0 -1.19040639897726e-05
Rx641 x641 0 1
Fxc641_640 x641 0 Vx640 -7.33991571995751
Cx641 x641 xm641 8.60345839298812e-13
Vx641 xm641 0 0
Gx641_1 x641 0 u1 0 8.73748264099121e-05
Rx642 x642 0 1
Fxc642_643 x642 0 Vx643 400.491826298254
Cx642 x642 xm642 9.68686303759719e-14
Vx642 xm642 0 0
Gx642_1 x642 0 u1 0 -3.44049552070881e-08
Rx643 x643 0 1
Fxc643_642 x643 0 Vx642 -1565.06631635724
Cx643 x643 xm643 9.68686303759719e-14
Vx643 xm643 0 0
Gx643_1 x643 0 u1 0 5.38460365103932e-05
Rx644 x644 0 1
Fxc644_645 x644 0 Vx645 42.1482081153883
Cx644 x644 xm644 1.48715507116435e-12
Vx644 xm644 0 0
Gx644_1 x644 0 u1 0 -7.86414618208791e-05
Rx645 x645 0 1
Fxc645_644 x645 0 Vx644 -67.5510389529967
Cx645 x645 xm645 1.48715507116435e-12
Vx645 xm645 0 0
Gx645_1 x645 0 u1 0 0.0053123124507828
Rx646 x646 0 1
Fxc646_647 x646 0 Vx647 146.063935401676
Cx646 x646 xm646 4.21127124032637e-13
Vx646 xm646 0 0
Gx646_1 x646 0 u1 0 -3.78915921294268e-07
Rx647 x647 0 1
Fxc647_646 x647 0 Vx646 -247.954240771237
Cx647 x647 xm647 4.21127124032637e-13
Vx647 xm647 0 0
Gx647_1 x647 0 u1 0 9.39538095806541e-05
Rx648 x648 0 1
Fxc648_649 x648 0 Vx649 582.017117759404
Cx648 x648 xm648 2.74413394468355e-13
Vx648 xm648 0 0
Gx648_1 x648 0 u1 0 -1.25127035678268e-07
Rx649 x649 0 1
Fxc649_648 x649 0 Vx648 -155.286726674999
Cx649 x649 xm649 2.74413394468355e-13
Vx649 xm649 0 0
Gx649_1 x649 0 u1 0 1.94305677890241e-05
Rx650 x650 0 1
Fxc650_651 x650 0 Vx651 60.3475739229705
Cx650 x650 xm650 1.53173944244712e-12
Vx650 xm650 0 0
Gx650_1 x650 0 u1 0 -1.64975116821098e-05
Rx651 x651 0 1
Fxc651_650 x651 0 Vx650 -51.0090617498541
Cx651 x651 xm651 1.53173944244712e-12
Vx651 xm651 0 0
Gx651_1 x651 0 u1 0 0.000841522592111678
Rx652 x652 0 1
Fxc652_653 x652 0 Vx653 80.9580092776718
Cx652 x652 xm652 1.91528411913751e-13
Vx652 xm652 0 0
Gx652_1 x652 0 u1 0 -1.36309480313815e-08
Rx653 x653 0 1
Fxc653_652 x653 0 Vx652 -2365.02486763484
Cx653 x653 xm653 1.91528411913751e-13
Vx653 xm653 0 0
Gx653_1 x653 0 u1 0 3.22375310636553e-05
Rx654 x654 0 1
Fxc654_655 x654 0 Vx655 5372.5869379414
Cx654 x654 xm654 2.36846187047956e-13
Vx654 xm654 0 0
Gx654_1 x654 0 u1 0 -7.64813940893495e-08
Rx655 x655 0 1
Fxc655_654 x655 0 Vx654 -28.0829381882011
Cx655 x655 xm655 2.36846187047956e-13
Vx655 xm655 0 0
Gx655_1 x655 0 u1 0 2.14782226275865e-06
Rx656 x656 0 1
Fxc656_657 x656 0 Vx657 19.3250670383103
Cx656 x656 xm656 8.29948243480383e-13
Vx656 xm656 0 0
Gx656_1 x656 0 u1 0 -3.57128851021728e-07
Rx657 x657 0 1
Fxc657_656 x657 0 Vx656 -576.762024552256
Cx657 x657 xm657 8.29948243480384e-13
Vx657 xm657 0 0
Gx657_1 x657 0 u1 0 0.000205978359141313
Rx658 x658 0 1
Fxc658_659 x658 0 Vx659 603.682156315705
Cx658 x658 xm658 1.49608073882079e-13
Vx658 xm658 0 0
Gx658_1 x658 0 u1 0 -3.29992362244313e-08
Rx659 x659 0 1
Fxc659_658 x659 0 Vx658 -543.970796589927
Cx659 x659 xm659 1.49608073882079e-13
Vx659 xm659 0 0
Gx659_1 x659 0 u1 0 1.79506208158631e-05
Rx660 x660 0 1
Fxc660_661 x660 0 Vx661 1322.1479610074
Cx660 x660 xm660 8.78155428912643e-14
Vx660 xm660 0 0
Gx660_1 x660 0 u1 0 -4.05492498989222e-09
Rx661 x661 0 1
Fxc661_660 x661 0 Vx660 -771.414078881183
Cx661 x661 xm661 8.78155428912643e-14
Vx661 xm661 0 0
Gx661_1 x661 0 u1 0 3.12802622601e-06
Rx662 x662 0 1
Fxc662_663 x662 0 Vx663 488.851824947172
Cx662 x662 xm662 4.67897291113138e-13
Vx662 xm662 0 0
Gx662_1 x662 0 u1 0 -1.16500297652523e-06
Rx663 x663 0 1
Fxc663_662 x663 0 Vx662 -57.7033107948782
Cx663 x663 xm663 4.67897291113138e-13
Vx663 xm663 0 0
Gx663_1 x663 0 u1 0 6.72245288313938e-05
Rx664 x664 0 1
Fxc664_665 x664 0 Vx665 151.888076613336
Cx664 x664 xm664 1.29257481425064e-13
Vx664 xm664 0 0
Gx664_1 x664 0 u1 0 -5.36857714448584e-09
Rx665 x665 0 1
Fxc665_664 x665 0 Vx664 -3231.7335928847
Cx665 x665 xm665 1.29257481425064e-13
Vx665 xm665 0 0
Gx665_1 x665 0 u1 0 1.73498111038279e-05
Rx666 x666 0 1
Fxc666_667 x666 0 Vx667 239.88755809339
Cx666 x666 xm666 1.14664608873347e-13
Vx666 xm666 0 0
Gx666_1 x666 0 u1 0 -2.93785468598374e-08
Rx667 x667 0 1
Fxc667_666 x667 0 Vx666 -1843.81500311164
Cx667 x667 xm667 1.14664608873347e-13
Vx667 xm667 0 0
Gx667_1 x667 0 u1 0 5.41686054697864e-05
Rx668 x668 0 1
Fxc668_669 x668 0 Vx669 70.9880716918783
Cx668 x668 xm668 1.69186391030051e-12
Vx668 xm668 0 0
Gx668_1 x668 0 u1 0 -1.0266195110642e-05
Rx669 x669 0 1
Fxc669_668 x669 0 Vx668 -45.3344820091232
Cx669 x669 xm669 1.69186391030051e-12
Vx669 xm669 0 0
Gx669_1 x669 0 u1 0 0.000465412637545548
Rx670 x670 0 1
Fxc670_671 x670 0 Vx671 73.6017611382118
Cx670 x670 xm670 5.92302008947924e-13
Vx670 xm670 0 0
Gx670_1 x670 0 u1 0 -2.2105564729806e-07
Rx671 x671 0 1
Fxc671_670 x671 0 Vx670 -364.965208422278
Cx671 x671 xm671 5.92302008947924e-13
Vx671 xm671 0 0
Gx671_1 x671 0 u1 0 8.0677620389058e-05
Rx672 x672 0 1
Fxc672_673 x672 0 Vx673 10.321898431088
Cx672 x672 xm672 1.69585389952454e-11
Vx672 xm672 0 0
Gx672_1 x672 0 u1 0 -0.0149627302145673
Rx673 x673 0 1
Fxc673_672 x673 0 Vx672 -4.18070048277477
Cx673 x673 xm673 1.69585389952454e-11
Vx673 xm673 0 0
Gx673_1 x673 0 u1 0 0.0625546934316702
Rx674 x674 0 1
Fxc674_675 x674 0 Vx675 27.859399188321
Cx674 x674 xm674 2.98300305540713e-12
Vx674 xm674 0 0
Gx674_1 x674 0 u1 0 -6.85669534759107e-05
Rx675 x675 0 1
Fxc675_674 x675 0 Vx674 -46.1111915730894
Cx675 x675 xm675 2.98300305540713e-12
Vx675 xm675 0 0
Gx675_1 x675 0 u1 0 0.00316170392731083
Rx676 x676 0 1
Fxc676_677 x676 0 Vx677 347.972586864213
Cx676 x676 xm676 1.26171155346877e-12
Vx676 xm676 0 0
Gx676_1 x676 0 u1 0 -4.02053090927509e-06
Rx677 x677 0 1
Fxc677_676 x677 0 Vx676 -18.0042127589785
Cx677 x677 xm677 1.26171155346877e-12
Vx677 xm677 0 0
Gx677_1 x677 0 u1 0 7.23864938946379e-05
Rx678 x678 0 1
Fxc678_679 x678 0 Vx679 1053.72686864721
Cx678 x678 xm678 2.40296590857126e-13
Vx678 xm678 0 0
Gx678_1 x678 0 u1 0 -9.56981518411347e-08
Rx679 x679 0 1
Fxc679_678 x679 0 Vx678 -175.312213273009
Cx679 x679 xm679 2.40296590857126e-13
Vx679 xm679 0 0
Gx679_1 x679 0 u1 0 1.67770548054058e-05
Rx680 x680 0 1
Fxc680_681 x680 0 Vx681 185.210931957782
Cx680 x680 xm680 7.07481712812474e-13
Vx680 xm680 0 0
Gx680_1 x680 0 u1 0 -7.95978269406673e-07
Rx681 x681 0 1
Fxc681_680 x681 0 Vx680 -117.683551508077
Cx681 x681 xm681 7.07481712812475e-13
Vx681 xm681 0 0
Gx681_1 x681 0 u1 0 9.36735496670306e-05
Rx682 x682 0 1
Fxc682_683 x682 0 Vx683 127.485127230105
Cx682 x682 xm682 2.47070341991198e-13
Vx682 xm682 0 0
Gx682_1 x682 0 u1 0 -1.78378091038833e-08
Rx683 x683 0 1
Fxc683_682 x683 0 Vx682 -1296.46356077898
Cx683 x683 xm683 2.47070341991198e-13
Vx683 xm683 0 0
Gx683_1 x683 0 u1 0 2.31260695073162e-05
Rx684 x684 0 1
Fxc684_685 x684 0 Vx685 3073.47289578065
Cx684 x684 xm684 6.42131520033378e-14
Vx684 xm684 0 0
Gx684_1 x684 0 u1 0 -5.01985648597099e-09
Rx685 x685 0 1
Fxc685_684 x685 0 Vx684 -715.518334451274
Cx685 x685 xm685 6.42131520033378e-14
Vx685 xm685 0 0
Gx685_1 x685 0 u1 0 3.59179935202639e-06
Rx686 x686 0 1
Fxc686_687 x686 0 Vx687 153.083418617645
Cx686 x686 xm686 1.12198183373626e-11
Vx686 xm686 0 0
Gx686_1 x686 0 u1 0 -0.00050521355718376
Rx687 x687 0 1
Fxc687_686 x687 0 Vx686 -1.11730418693402
Cx687 x687 xm687 1.12198183373626e-11
Vx687 xm687 0 0
Gx687_1 x687 0 u1 0 0.000564477222737245
Rx688 x688 0 1
Fxc688_689 x688 0 Vx689 4.46659079740919
Cx688 x688 xm688 3.2472763080511e-12
Vx688 xm688 0 0
Gx688_1 x688 0 u1 0 -1.92382673676807e-05
Rx689 x689 0 1
Fxc689_688 x689 0 Vx688 -257.732822465335
Cx689 x689 xm689 3.2472763080511e-12
Vx689 xm689 0 0
Gx689_1 x689 0 u1 0 0.00495833294801508
Rx690 x690 0 1
Fxc690_691 x690 0 Vx691 0.920155029332168
Cx690 x690 xm690 3.71285809172693e-12
Vx690 xm690 0 0
Gx690_1 x690 0 u1 0 -2.52299541872688e-06
Rx691 x691 0 1
Fxc691_690 x691 0 Vx690 -1047.88094678809
Cx691 x691 xm691 3.71285809172693e-12
Vx691 xm691 0 0
Gx691_1 x691 0 u1 0 0.00264379882811754
Rx692 x692 0 1
Fxc692_693 x692 0 Vx693 28.4620874667522
Cx692 x692 xm692 7.59177081056463e-13
Vx692 xm692 0 0
Gx692_1 x692 0 u1 0 -1.34912766447843e-07
Rx693 x693 0 1
Fxc693_692 x693 0 Vx692 -778.086552589465
Cx693 x693 xm693 7.59177081056463e-13
Vx693 xm693 0 0
Gx693_1 x693 0 u1 0 0.00010497380934571
Rx694 x694 0 1
Fxc694_695 x694 0 Vx695 93.0505482090238
Cx694 x694 xm694 2.02585528546519e-13
Vx694 xm694 0 0
Gx694_1 x694 0 u1 0 -1.05325412110591e-08
Rx695 x695 0 1
Fxc695_694 x695 0 Vx694 -3204.2871633725
Cx695 x695 xm695 2.02585528546519e-13
Vx695 xm695 0 0
Gx695_1 x695 0 u1 0 3.37492866002886e-05
Rx696 x696 0 1
Fxc696_697 x696 0 Vx697 3843.42632853417
Cx696 x696 xm696 4.24372223574733e-14
Vx696 xm696 0 0
Gx696_1 x696 0 u1 0 -3.67750135030707e-09
Rx697 x697 0 1
Fxc697_696 x697 0 Vx696 -1963.13659128213
Cx697 x697 xm697 4.24372223574733e-14
Vx697 xm697 0 0
Gx697_1 x697 0 u1 0 7.21943746527724e-06
Rx698 x698 0 1
Fxc698_699 x698 0 Vx699 38139.7686075898
Cx698 x698 xm698 1.00885100580125e-13
Vx698 xm698 0 0
Gx698_1 x698 0 u1 0 -1.84351238854034e-08
Rx699 x699 0 1
Fxc699_698 x699 0 Vx698 -37.6313475280237
Cx699 x699 xm699 1.00885100580125e-13
Vx699 xm699 0 0
Gx699_1 x699 0 u1 0 6.93738553653786e-07
Rx700 x700 0 1
Fxc700_701 x700 0 Vx701 254.641692644996
Cx700 x700 xm700 4.00195036079336e-13
Vx700 xm700 0 0
Gx700_1 x700 0 u1 0 -1.25786388027372e-07
Rx701 x701 0 1
Fxc701_700 x701 0 Vx700 -286.045823131594
Cx701 x701 xm701 4.00195036079336e-13
Vx701 xm701 0 0
Gx701_1 x701 0 u1 0 3.59806709020398e-05
Rx702 x702 0 1
Fxc702_703 x702 0 Vx703 275.460269286693
Cx702 x702 xm702 2.78329702880848e-13
Vx702 xm702 0 0
Gx702_1 x702 0 u1 0 -1.55192192330146e-08
Rx703 x703 0 1
Fxc703_702 x703 0 Vx702 -712.188250368702
Cx703 x703 xm703 2.78329702880848e-13
Vx703 xm703 0 0
Gx703_1 x703 0 u1 0 1.1052605592649e-05
Rx704 x704 0 1
Fxc704_705 x704 0 Vx705 54.089280062518
Cx704 x704 xm704 1.59370707888504e-12
Vx704 xm704 0 0
Gx704_1 x704 0 u1 0 -3.41145821417576e-06
Rx705 x705 0 1
Fxc705_704 x705 0 Vx704 -122.453170282091
Cx705 x705 xm705 1.59370707888504e-12
Vx705 xm705 0 0
Gx705_1 x705 0 u1 0 0.000417743873610703
Rx706 x706 0 1
Fxc706_707 x706 0 Vx707 245.077982928638
Cx706 x706 xm706 1.50328460311422e-12
Vx706 xm706 0 0
Gx706_1 x706 0 u1 0 -4.47339931597085e-06
Rx707 x707 0 1
Fxc707_706 x707 0 Vx706 -32.0446757856762
Cx707 x707 xm707 1.50328460311422e-12
Vx707 xm707 0 0
Gx707_1 x707 0 u1 0 0.000143348630740151
Rx708 x708 0 1
Fxc708_709 x708 0 Vx709 122.306784606395
Cx708 x708 xm708 2.99713440633919e-12
Vx708 xm708 0 0
Gx708_1 x708 0 u1 0 -3.80802278572733e-05
Rx709 x709 0 1
Fxc709_708 x709 0 Vx708 -15.0224505795789
Cx709 x709 xm709 2.99713440633919e-12
Vx709 xm709 0 0
Gx709_1 x709 0 u1 0 0.000572058341044993
Rx710 x710 0 1
Fxc710_711 x710 0 Vx711 325.182194033925
Cx710 x710 xm710 4.59729955117924e-13
Vx710 xm710 0 0
Gx710_1 x710 0 u1 0 -6.99533686796408e-08
Rx711 x711 0 1
Fxc711_710 x711 0 Vx710 -229.506743200215
Cx711 x711 xm711 4.59729955117924e-13
Vx711 xm711 0 0
Gx711_1 x711 0 u1 0 1.60547698215483e-05
Rx712 x712 0 1
Fxc712_713 x712 0 Vx713 6.65135965755537
Cx712 x712 xm712 2.42031501813512e-12
Vx712 xm712 0 0
Gx712_1 x712 0 u1 0 -2.00800784133623e-06
Rx713 x713 0 1
Fxc713_712 x713 0 Vx712 -466.419665326437
Cx713 x713 xm713 2.42031501813512e-12
Vx713 xm713 0 0
Gx713_1 x713 0 u1 0 0.000936574345328907
Rx714 x714 0 1
Fxc714_715 x714 0 Vx715 1.09594520754942
Cx714 x714 xm714 5.54877528405509e-13
Vx714 xm714 0 0
Gx714_1 x714 0 u1 0 -7.58034550626094e-10
Rx715 x715 0 1
Fxc715_714 x715 0 Vx714 -56822.6373554408
Cx715 x715 xm715 5.54877528405509e-13
Vx715 xm715 0 0
Gx715_1 x715 0 u1 0 4.30735223731211e-05
Rx716 x716 0 1
Cx716 x716 0 1.61089900076846e-09
Gx716_1 x716 0 u1 0 -0.380021832809238
Rx717 x717 0 1
Fxc717_718 x717 0 Vx718 0.983027769254327
Cx717 x717 xm717 2.19812424587013e-10
Vx717 xm717 0 0
Gx717_1 x717 0 u1 0 -0.0164369770428683
Rx718 x718 0 1
Fxc718_717 x718 0 Vx717 -8.61137872719285
Cx718 x718 xm718 2.19812424587013e-10
Vx718 xm718 0 0
Gx718_1 x718 0 u1 0 0.141545034446313
Rx719 x719 0 1
Fxc719_720 x719 0 Vx720 9.23069240641804
Cx719 x719 xm719 1.87705184078918e-09
Vx719 xm719 0 0
Gx719_1 x719 0 u1 0 -0.074486287007802
Rx720 x720 0 1
Fxc720_719 x720 0 Vx719 -0.132068389727408
Cx720 x720 xm720 1.87705184078918e-09
Vx720 xm720 0 0
Gx720_1 x720 0 u1 0 0.00983728398189393
Rx721 x721 0 1
Fxc721_722 x721 0 Vx722 7.61541940666506
Cx721 x721 xm721 4.32510417049148e-11
Vx721 xm721 0 0
Gx721_1 x721 0 u1 0 -1.71438375362709e-06
Rx722 x722 0 1
Fxc722_721 x722 0 Vx721 -158.123974658734
Cx722 x722 xm722 4.32510417049148e-11
Vx722 xm722 0 0
Gx722_1 x722 0 u1 0 0.000271085173213875
Rx723 x723 0 1
Fxc723_724 x723 0 Vx724 223.966016863591
Cx723 x723 xm723 6.12250410889856e-12
Vx723 xm723 0 0
Gx723_1 x723 0 u1 0 -7.33981667417477e-07
Rx724 x724 0 1
Fxc724_723 x724 0 Vx723 -131.544849629263
Cx724 x724 xm724 6.12250410889856e-12
Vx724 xm724 0 0
Gx724_1 x724 0 u1 0 9.6551508071068e-05
Rx725 x725 0 1
Fxc725_726 x725 0 Vx726 454.493702970474
Cx725 x725 xm725 4.14799482577559e-11
Vx725 xm725 0 0
Gx725_1 x725 0 u1 0 -0.00666731448011287
Rx726 x726 0 1
Fxc726_725 x726 0 Vx725 -0.0697268883519739
Cx726 x726 xm726 4.14799482577559e-11
Vx726 xm726 0 0
Gx726_1 x726 0 u1 0 0.000464891092362329
Rx727 x727 0 1
Fxc727_728 x727 0 Vx728 4036.97442282991
Cx727 x727 xm727 1.45549226115441e-14
Vx727 xm727 0 0
Gx727_1 x727 0 u1 0 -2.06700273833501e-10
Rx728 x728 0 1
Fxc728_727 x728 0 Vx727 -24028.3143574083
Cx728 x728 xm728 1.45549226115441e-14
Vx728 xm728 0 0
Gx728_1 x728 0 u1 0 4.96665915743375e-06
Rx729 x729 0 1
Fxc729_730 x729 0 Vx730 17.3301584740127
Cx729 x729 xm729 1.60409482204103e-11
Vx729 xm729 0 0
Gx729_1 x729 0 u1 0 -0.000508184969198248
Rx730 x730 0 1
Fxc730_729 x730 0 Vx729 -8.00923470638368
Cx730 x730 xm730 1.60409482204104e-11
Vx730 xm730 0 0
Gx730_1 x730 0 u1 0 0.00407017269256513
Rx731 x731 0 1
Fxc731_732 x731 0 Vx732 5.02306883287156
Cx731 x731 xm731 1.87789127101595e-11
Vx731 xm731 0 0
Gx731_1 x731 0 u1 0 -0.000141186579965918
Rx732 x732 0 1
Fxc732_731 x732 0 Vx731 -43.1965037584085
Cx732 x732 xm732 1.87789127101595e-11
Vx732 xm732 0 0
Gx732_1 x732 0 u1 0 0.00609876663213461
Rx733 x733 0 1
Fxc733_734 x733 0 Vx734 90.9668866205123
Cx733 x733 xm733 1.4701859252872e-12
Vx733 xm733 0 0
Gx733_1 x733 0 u1 0 -6.01294552206778e-07
Rx734 x734 0 1
Fxc734_733 x734 0 Vx733 -133.79088771572
Cx734 x734 xm734 1.4701859252872e-12
Vx734 xm734 0 0
Gx734_1 x734 0 u1 0 8.04477319183712e-05
Rx735 x735 0 1
Fxc735_736 x735 0 Vx736 41.8858479213457
Cx735 x735 xm735 2.39937551270491e-13
Vx735 xm735 0 0
Gx735_1 x735 0 u1 0 -1.53317648104001e-09
Rx736 x736 0 1
Fxc736_735 x736 0 Vx735 -9338.99859179738
Cx736 x736 xm736 2.39937551270491e-13
Vx736 xm736 0 0
Gx736_1 x736 0 u1 0 1.43183329974096e-05
Rx737 x737 0 1
Fxc737_738 x737 0 Vx738 1716.10105074822
Cx737 x737 xm737 3.58178612159909e-13
Vx737 xm737 0 0
Gx737_1 x737 0 u1 0 -2.92729758772931e-08
Rx738 x738 0 1
Fxc738_737 x738 0 Vx737 -124.757891915171
Cx738 x738 xm738 3.58178612159909e-13
Vx738 xm738 0 0
Gx738_1 x738 0 u1 0 3.65203476053475e-06
Rx739 x739 0 1
Fxc739_740 x739 0 Vx740 45.2313098936706
Cx739 x739 xm739 5.21591991919758e-12
Vx739 xm739 0 0
Gx739_1 x739 0 u1 0 -1.78805384035417e-05
Rx740 x740 0 1
Fxc740_739 x740 0 Vx739 -58.4192728832078
Cx740 x740 xm740 5.21591991919758e-12
Vx740 xm740 0 0
Gx740_1 x740 0 u1 0 0.00104456805229518
Rx741 x741 0 1
Fxc741_742 x741 0 Vx742 8.1505522628012
Cx741 x741 xm741 9.36281020722464e-13
Vx741 xm741 0 0
Gx741_1 x741 0 u1 0 -2.50435299111019e-08
Rx742 x742 0 1
Fxc742_741 x742 0 Vx741 -3313.29304439357
Cx742 x742 xm742 9.36281020722465e-13
Vx742 xm742 0 0
Gx742_1 x742 0 u1 0 8.29765534615162e-05
Rx743 x743 0 1
Fxc743_744 x743 0 Vx744 325.027711282142
Cx743 x743 xm743 5.00909331659054e-13
Vx743 xm743 0 0
Gx743_1 x743 0 u1 0 -1.13988359722108e-08
Rx744 x744 0 1
Fxc744_743 x744 0 Vx743 -742.362475278835
Cx744 x744 xm744 5.00909331659054e-13
Vx744 xm744 0 0
Gx744_1 x744 0 u1 0 8.46206808762783e-06
Rx745 x745 0 1
Fxc745_746 x745 0 Vx746 576.655639001651
Cx745 x745 xm745 2.21603934379445e-12
Vx745 xm745 0 0
Gx745_1 x745 0 u1 0 -1.14731910751247e-06
Rx746 x746 0 1
Fxc746_745 x746 0 Vx745 -16.9723903845247
Cx746 x746 xm746 2.21603934379445e-12
Vx746 xm746 0 0
Gx746_1 x746 0 u1 0 1.94727477883261e-05
Rx747 x747 0 1
Fxc747_748 x747 0 Vx748 266596.978331078
Cx747 x747 xm747 1.03257318571619e-14
Vx747 xm747 0 0
Gx747_1 x747 0 u1 0 -1.32187256858776e-09
Rx748 x748 0 1
Fxc748_747 x748 0 Vx747 -1162.75242451968
Cx748 x748 xm748 1.03257318571619e-14
Vx748 xm748 0 0
Gx748_1 x748 0 u1 0 1.53701053403147e-06
Rx749 x749 0 1
Fxc749_750 x749 0 Vx750 2252.24869682317
Cx749 x749 xm749 2.74819843338129e-12
Vx749 xm749 0 0
Gx749_1 x749 0 u1 0 -6.85233013483777e-06
Rx750 x750 0 1
Fxc750_749 x750 0 Vx749 -1.77478002706601
Cx750 x750 xm750 2.74819843338129e-12
Vx750 xm750 0 0
Gx750_1 x750 0 u1 0 1.21613786621726e-05
Rx751 x751 0 1
Fxc751_752 x751 0 Vx752 569.330456169478
Cx751 x751 xm751 4.24036342517206e-12
Vx751 xm751 0 0
Gx751_1 x751 0 u1 0 -6.87874744809385e-06
Rx752 x752 0 1
Fxc752_751 x752 0 Vx751 -4.3657164348973
Cx752 x752 xm752 4.24036342517206e-12
Vx752 xm752 0 0
Gx752_1 x752 0 u1 0 3.00306607856512e-05
Rx753 x753 0 1
Fxc753_754 x753 0 Vx754 550.949593871042
Cx753 x753 xm753 9.58496587203372e-13
Vx753 xm753 0 0
Gx753_1 x753 0 u1 0 -2.10785269545362e-07
Rx754 x754 0 1
Fxc754_753 x754 0 Vx753 -82.1982470199113
Cx754 x754 xm754 9.58496587203372e-13
Vx754 xm754 0 0
Gx754_1 x754 0 u1 0 1.73261796542482e-05
Rx755 x755 0 1
Fxc755_756 x755 0 Vx756 182.97171001156
Cx755 x755 xm755 1.12815467078128e-12
Vx755 xm755 0 0
Gx755_1 x755 0 u1 0 -2.37610595248639e-07
Rx756 x756 0 1
Fxc756_755 x756 0 Vx755 -153.792395896455
Cx756 x756 xm756 1.12815467078128e-12
Vx756 xm756 0 0
Gx756_1 x756 0 u1 0 3.65427027336711e-05
Rx757 x757 0 1
Fxc757_758 x757 0 Vx758 37.5576872473799
Cx757 x757 xm757 1.79517864865178e-12
Vx757 xm757 0 0
Gx757_1 x757 0 u1 0 -8.02933638059489e-07
Rx758 x758 0 1
Fxc758_757 x758 0 Vx757 -254.619351087646
Cx758 x758 xm758 1.79517864865178e-12
Vx758 xm758 0 0
Gx758_1 x758 0 u1 0 0.00020444244188915
Rx759 x759 0 1
Fxc759_760 x759 0 Vx760 855.826912858585
Cx759 x759 xm759 6.11941306890275e-13
Vx759 xm759 0 0
Gx759_1 x759 0 u1 0 -1.63648126752286e-07
Rx760 x760 0 1
Fxc760_759 x760 0 Vx759 -72.4651464577562
Cx760 x760 xm760 6.11941306890275e-13
Vx760 xm760 0 0
Gx760_1 x760 0 u1 0 1.18587854726419e-05
Rx761 x761 0 1
Fxc761_762 x761 0 Vx762 31.0114861002044
Cx761 x761 xm761 1.42015889054634e-12
Vx761 xm761 0 0
Gx761_1 x761 0 u1 0 -6.60416903333314e-08
Rx762 x762 0 1
Fxc762_761 x762 0 Vx761 -853.233536461557
Cx762 x762 xm762 1.42015889054634e-12
Vx762 xm762 0 0
Gx762_1 x762 0 u1 0 5.63489849970073e-05
Rx763 x763 0 1
Fxc763_764 x763 0 Vx764 39.4045000736137
Cx763 x763 xm763 7.91863406834521e-12
Vx763 xm763 0 0
Gx763_1 x763 0 u1 0 -7.79911380437587e-05
Rx764 x764 0 1
Fxc764_763 x764 0 Vx763 -29.0405149593984
Cx764 x764 xm764 7.91863406834521e-12
Vx764 xm764 0 0
Gx764_1 x764 0 u1 0 0.00226490281106028
Rx765 x765 0 1
Fxc765_766 x765 0 Vx766 1550.50038070534
Cx765 x765 xm765 9.12011682999143e-13
Vx765 xm765 0 0
Gx765_1 x765 0 u1 0 -6.89597511019354e-08
Rx766 x766 0 1
Fxc766_765 x766 0 Vx765 -65.5514663246482
Cx766 x766 xm766 9.12011682999143e-13
Vx766 xm766 0 0
Gx766_1 x766 0 u1 0 4.52041280211464e-06
Rx767 x767 0 1
Fxc767_768 x767 0 Vx768 131.98632194045
Cx767 x767 xm767 2.64454642404486e-12
Vx767 xm767 0 0
Gx767_1 x767 0 u1 0 -4.06385100249608e-07
Rx768 x768 0 1
Fxc768_767 x768 0 Vx767 -101.366474128854
Cx768 x768 xm768 2.64454642404486e-12
Vx768 xm768 0 0
Gx768_1 x768 0 u1 0 4.11938247508035e-05
Rx769 x769 0 1
Fxc769_770 x769 0 Vx770 31.5118028228
Cx769 x769 xm769 1.51286572624691e-11
Vx769 xm769 0 0
Gx769_1 x769 0 u1 0 -4.32140540469364e-05
Rx770 x770 0 1
Fxc770_769 x770 0 Vx769 -18.6443156098518
Cx770 x770 xm770 1.51286572624691e-11
Vx770 xm770 0 0
Gx770_1 x770 0 u1 0 0.000805696462432276
Rx771 x771 0 1
Fxc771_772 x771 0 Vx772 4.17455736131485
Cx771 x771 xm771 1.22419165937248e-10
Vx771 xm771 0 0
Gx771_1 x771 0 u1 0 -0.00957186809740095
Rx772 x772 0 1
Fxc772_771 x772 0 Vx771 -5.03704227937591
Cx772 x772 xm772 1.22419165937248e-10
Vx772 xm772 0 0
Gx772_1 x772 0 u1 0 0.0482139042992181
Rx773 x773 0 1
Fxc773_774 x773 0 Vx774 109.634258986536
Cx773 x773 xm773 1.76967136661136e-11
Vx773 xm773 0 0
Gx773_1 x773 0 u1 0 -2.46339135708522e-05
Rx774 x774 0 1
Fxc774_773 x774 0 Vx773 -6.18998837559069
Cx774 x774 xm774 1.76967136661136e-11
Vx774 xm774 0 0
Gx774_1 x774 0 u1 0 0.000152483638648881
Rx775 x775 0 1
Fxc775_776 x775 0 Vx776 1.11486755016664
Cx775 x775 xm775 1.26800162802138e-11
Vx775 xm775 0 0
Gx775_1 x775 0 u1 0 -2.11716806993752e-07
Rx776 x776 0 1
Fxc776_775 x776 0 Vx775 -1435.83336212759
Cx776 x776 xm776 1.26800162802138e-11
Vx776 xm776 0 0
Gx776_1 x776 0 u1 0 0.000303990054804757
Rx777 x777 0 1
Cx777 x777 0 7.05227504597919e-09
Gx777_1 x777 0 u1 0 -0.372335092042141
Rx778 x778 0 1
Fxc778_779 x778 0 Vx779 240.422659858283
Cx778 x778 xm778 1.15460286288366e-12
Vx778 xm778 0 0
Gx778_1 x778 0 u1 0 -2.27633662567822e-07
Rx779 x779 0 1
Fxc779_778 x779 0 Vx778 -119.781114034112
Cx779 x779 xm779 1.15460286288366e-12
Vx779 xm779 0 0
Gx779_1 x779 0 u1 0 2.72662136940388e-05
Rx780 x780 0 1
Fxc780_781 x780 0 Vx781 3.29276953715306
Cx780 x780 xm780 2.18132271178657e-10
Vx780 xm780 0 0
Gx780_1 x780 0 u1 0 -9.01818336091932e-06
Rx781 x781 0 1
Fxc781_780 x781 0 Vx780 -98.2011932925076
Cx781 x781 xm781 2.18132271178657e-10
Vx781 xm781 0 0
Gx781_1 x781 0 u1 0 0.000885596367372914
Rx782 x782 0 1
Fxc782_783 x782 0 Vx783 8.21682672361746
Cx782 x782 xm782 8.40037698819289e-11
Vx782 xm782 0 0
Gx782_1 x782 0 u1 0 -0.00116952752666867
Rx783 x783 0 1
Fxc783_782 x783 0 Vx782 -8.06037132510542
Cx783 x783 xm783 8.40037698819289e-11
Vx783 xm783 0 0
Gx783_1 x783 0 u1 0 0.00942682613988161
Rx784 x784 0 1
Fxc784_785 x784 0 Vx785 5.7526568772806
Cx784 x784 xm784 5.30998399535694e-11
Vx784 xm784 0 0
Gx784_1 x784 0 u1 0 -2.55299070295937e-05
Rx785 x785 0 1
Fxc785_784 x785 0 Vx784 -42.5986970334547
Cx785 x785 xm785 5.30998399535694e-11
Vx785 xm785 0 0
Gx785_1 x785 0 u1 0 0.00108754077484593
Rx786 x786 0 1
Fxc786_787 x786 0 Vx787 535.33343695727
Cx786 x786 xm786 1.35912169198298e-12
Vx786 xm786 0 0
Gx786_1 x786 0 u1 0 -1.3480326242589e-07
Rx787 x787 0 1
Fxc787_786 x787 0 Vx786 -102.630190274221
Cx787 x787 xm787 1.35912169198298e-12
Vx787 xm787 0 0
Gx787_1 x787 0 u1 0 1.38348844723548e-05
Rx788 x788 0 1
Fxc788_789 x788 0 Vx789 47.105537377694
Cx788 x788 xm788 6.31264225400471e-12
Vx788 xm788 0 0
Gx788_1 x788 0 u1 0 -2.90961458202697e-06
Rx789 x789 0 1
Fxc789_788 x789 0 Vx788 -58.5677360242781
Cx789 x789 xm789 6.31264225400471e-12
Vx789 xm789 0 0
Gx789_1 x789 0 u1 0 0.000170409538772546
Rx790 x790 0 1
Fxc790_791 x790 0 Vx791 0.720801659391959
Cx790 x790 xm790 1.33436643953763e-11
Vx790 xm790 0 0
Gx790_1 x790 0 u1 0 -1.4135923694065e-06
Rx791 x791 0 1
Fxc791_790 x791 0 Vx790 -1159.83401597914
Cx791 x791 xm791 1.33436643953763e-11
Vx791 xm791 0 0
Gx791_1 x791 0 u1 0 0.00163953251476621
Rx792 x792 0 1
Fxc792_793 x792 0 Vx793 443.928905607266
Cx792 x792 xm792 1.32642627349223e-11
Vx792 xm792 0 0
Gx792_1 x792 0 u1 0 -6.69400185299945e-06
Rx793 x793 0 1
Fxc793_792 x793 0 Vx792 -3.9409703838887
Cx793 x793 xm793 1.32642627349223e-11
Vx793 xm793 0 0
Gx793_1 x793 0 u1 0 2.63808630523669e-05
Rx794 x794 0 1
Fxc794_795 x794 0 Vx795 23.8032819070874
Cx794 x794 xm794 1.08698420955425e-11
Vx794 xm794 0 0
Gx794_1 x794 0 u1 0 -5.024048330275e-06
Rx795 x795 0 1
Fxc795_794 x795 0 Vx794 -63.0733320089588
Cx795 x795 xm795 1.08698420955425e-11
Vx795 xm795 0 0
Gx795_1 x795 0 u1 0 0.00031688346836449
Rx796 x796 0 1
Fxc796_797 x796 0 Vx797 97.250099169652
Cx796 x796 xm796 4.56998680318091e-12
Vx796 xm796 0 0
Gx796_1 x796 0 u1 0 -2.05887946944537e-06
Rx797 x797 0 1
Fxc797_796 x797 0 Vx796 -75.2886756000796
Cx797 x797 xm797 4.56998680318091e-12
Vx797 xm797 0 0
Gx797_1 x797 0 u1 0 0.000155010308474736
Rx798 x798 0 1
Cx798 x798 0 1.02081938428761e-08
Gx798_1 x798 0 u1 0 -0.273298145902074
Rx799 x799 0 1
Fxc799_800 x799 0 Vx800 14.3639677855823
Cx799 x799 xm799 1.53254609092949e-11
Vx799 xm799 0 0
Gx799_1 x799 0 u1 0 -2.75211978087786e-06
Rx800 x800 0 1
Fxc800_799 x800 0 Vx799 -126.887548866497
Cx800 x800 xm800 1.53254609092949e-11
Vx800 xm800 0 0
Gx800_1 x800 0 u1 0 0.000349209733182593
Rx801 x801 0 1
Cx801 x801 0 5.04506053260489e-08
Gx801_1 x801 0 u1 0 -0.237497172545955
Rx802 x802 0 1
Cx802 x802 0 3.53627063161835e-13
Gx802_2 x802 0 u2 0 -78.4311936160815
Rx803 x803 0 1
Cx803 x803 0 8.59855014759414e-12
Gx803_2 x803 0 u2 0 -490.320531339327
Rx804 x804 0 1
Fxc804_805 x804 0 Vx805 111.946950651084
Cx804 x804 xm804 1.52013265599724e-13
Vx804 xm804 0 0
Gx804_2 x804 0 u2 0 -0.0448639665961424
Rx805 x805 0 1
Fxc805_804 x805 0 Vx804 -73.0620408934091
Cx805 x805 xm805 1.52013265599724e-13
Vx805 xm805 0 0
Gx805_2 x805 0 u2 0 3.27785296208789
Rx806 x806 0 1
Fxc806_807 x806 0 Vx807 78.1460349279812
Cx806 x806 xm806 1.34030288980988e-11
Vx806 xm806 0 0
Gx806_2 x806 0 u2 0 -418.395448073798
Rx807 x807 0 1
Fxc807_806 x807 0 Vx806 -0.00756161147043389
Cx807 x807 xm807 1.34030288980988e-11
Vx807 xm807 0 0
Gx807_2 x807 0 u2 0 3.16374381933216
Rx808 x808 0 1
Fxc808_809 x808 0 Vx809 560.182600379328
Cx808 x808 xm808 3.10934658884836e-14
Vx808 xm808 0 0
Gx808_2 x808 0 u2 0 -9.11988505452926e-07
Rx809 x809 0 1
Fxc809_808 x809 0 Vx808 -469.469560608369
Cx809 x809 xm809 3.10934658884836e-14
Vx809 xm809 0 0
Gx809_2 x809 0 u2 0 0.000428150842934869
Rx810 x810 0 1
Fxc810_811 x810 0 Vx811 21467.4775020896
Cx810 x810 xm810 8.40733664871429e-15
Vx810 xm810 0 0
Gx810_2 x810 0 u2 0 -4.61440373837623e-08
Rx811 x811 0 1
Fxc811_810 x811 0 Vx810 -169.230255222059
Cx811 x811 xm811 8.40733664871429e-15
Vx811 xm811 0 0
Gx811_2 x811 0 u2 0 7.80896722343033e-06
Rx812 x812 0 1
Fxc812_813 x812 0 Vx813 17279.2782798773
Cx812 x812 xm812 1.94523784543502e-15
Vx812 xm812 0 0
Gx812_2 x812 0 u2 0 -1.13957347418057e-09
Rx813 x813 0 1
Fxc813_812 x813 0 Vx812 -3945.09077931237
Cx813 x813 xm813 1.94523784543502e-15
Vx813 xm813 0 0
Gx813_2 x813 0 u2 0 4.49572080533873e-06
Rx814 x814 0 1
Fxc814_815 x814 0 Vx815 534.100178275924
Cx814 x814 xm814 1.91730724654873e-14
Vx814 xm814 0 0
Gx814_2 x814 0 u2 0 -1.31971590144073e-07
Rx815 x815 0 1
Fxc815_814 x815 0 Vx814 -1322.64424794249
Cx815 x815 xm815 1.91730724654873e-14
Vx815 xm815 0 0
Gx815_2 x815 0 u2 0 0.000174551464595882
Rx816 x816 0 1
Fxc816_817 x816 0 Vx817 51.0602372944747
Cx816 x816 xm816 4.56584091846018e-14
Vx816 xm816 0 0
Gx816_2 x816 0 u2 0 -3.45972745266959e-07
Rx817 x817 0 1
Fxc817_816 x817 0 Vx816 -2454.7487115417
Cx817 x817 xm817 4.56584091846018e-14
Vx817 xm817 0 0
Gx817_2 x817 0 u2 0 0.000849276150672613
Rx818 x818 0 1
Fxc818_819 x818 0 Vx819 550120.787252286
Cx818 x818 xm818 6.22970485029519e-16
Vx818 xm818 0 0
Gx818_2 x818 0 u2 0 -3.0547376018853e-10
Rx819 x819 0 1
Fxc819_818 x819 0 Vx818 -1229.74008330112
Cx819 x819 xm819 6.22970485029519e-16
Vx819 xm819 0 0
Gx819_2 x819 0 u2 0 3.7565332730055e-07
Rx820 x820 0 1
Fxc820_821 x820 0 Vx821 12.7664587590957
Cx820 x820 xm820 1.1019165711965e-12
Vx820 xm820 0 0
Gx820_2 x820 0 u2 0 -0.160546600712626
Rx821 x821 0 1
Fxc821_820 x821 0 Vx820 -18.7364216141508
Cx821 x821 xm821 1.1019165711965e-12
Vx821 xm821 0 0
Gx821_2 x821 0 u2 0 3.00806879967048
Rx822 x822 0 1
Fxc822_823 x822 0 Vx823 15258.1856472676
Cx822 x822 xm822 4.28178588649374e-16
Vx822 xm822 0 0
Gx822_2 x822 0 u2 0 -2.69993939959885e-10
Rx823 x823 0 1
Fxc823_822 x823 0 Vx822 -94575.535325067
Cx823 x823 xm823 4.28178588649374e-16
Vx823 xm823 0 0
Gx823_2 x823 0 u2 0 2.55348214062302e-05
Rx824 x824 0 1
Fxc824_825 x824 0 Vx825 7780.24516947265
Cx824 x824 xm824 2.43387977270851e-14
Vx824 xm824 0 0
Gx824_2 x824 0 u2 0 -3.93387593242905e-07
Rx825 x825 0 1
Fxc825_824 x825 0 Vx824 -57.5833395090103
Cx825 x825 xm825 2.43387977270851e-14
Vx825 xm825 0 0
Gx825_2 x825 0 u2 0 2.26525713403386e-05
Rx826 x826 0 1
Fxc826_827 x826 0 Vx827 156.713786566692
Cx826 x826 xm826 1.05011663800036e-13
Vx826 xm826 0 0
Gx826_2 x826 0 u2 0 -2.26427023507671e-05
Rx827 x827 0 1
Fxc827_826 x827 0 Vx826 -154.802365874463
Cx827 x827 xm827 1.05011663800036e-13
Vx827 xm827 0 0
Gx827_2 x827 0 u2 0 0.00350514389369
Rx828 x828 0 1
Fxc828_829 x828 0 Vx829 390.683198738113
Cx828 x828 xm828 1.08883637079586e-14
Vx828 xm828 0 0
Gx828_2 x828 0 u2 0 -1.19957849738671e-08
Rx829 x829 0 1
Fxc829_828 x829 0 Vx828 -5816.91372281582
Cx829 x829 xm829 1.08883637079586e-14
Vx829 xm829 0 0
Gx829_2 x829 0 u2 0 6.97784462304354e-05
Rx830 x830 0 1
Fxc830_831 x830 0 Vx831 1041.13125074382
Cx830 x830 xm830 1.79569174984714e-14
Vx830 xm830 0 0
Gx830_2 x830 0 u2 0 -1.46900605498445e-07
Rx831 x831 0 1
Fxc831_830 x831 0 Vx830 -806.957748296937
Cx831 x831 xm831 1.79569174984714e-14
Vx831 xm831 0 0
Gx831_2 x831 0 u2 0 0.000118542581836482
Rx832 x832 0 1
Fxc832_833 x832 0 Vx833 1057.0564537887
Cx832 x832 xm832 1.89102617067545e-14
Vx832 xm832 0 0
Gx832_2 x832 0 u2 0 -1.61268368869956e-07
Rx833 x833 0 1
Fxc833_832 x833 0 Vx832 -720.302576869593
Cx833 x833 xm833 1.89102617067545e-14
Vx833 xm833 0 0
Gx833_2 x833 0 u2 0 0.000116162021664585
Rx834 x834 0 1
Fxc834_835 x834 0 Vx835 7156.78813973339
Cx834 x834 xm834 1.08306461059872e-14
Vx834 xm834 0 0
Gx834_2 x834 0 u2 0 -4.38716048950967e-08
Rx835 x835 0 1
Fxc835_834 x835 0 Vx834 -326.12687828736
Cx835 x835 xm835 1.08306461059872e-14
Vx835 xm835 0 0
Gx835_2 x835 0 u2 0 1.43077095498943e-05
Rx836 x836 0 1
Fxc836_837 x836 0 Vx837 13.646492462318
Cx836 x836 xm836 2.09659001892218e-13
Vx836 xm836 0 0
Gx836_2 x836 0 u2 0 -0.000168504476669207
Rx837 x837 0 1
Fxc837_836 x837 0 Vx836 -467.327802517942
Cx837 x837 xm837 2.09659001892218e-13
Vx837 xm837 0 0
Gx837_2 x837 0 u2 0 0.0787468267962561
Rx838 x838 0 1
Fxc838_839 x838 0 Vx839 2415.37622901448
Cx838 x838 xm838 1.6602740464064e-14
Vx838 xm838 0 0
Gx838_2 x838 0 u2 0 -8.34054652355412e-08
Rx839 x839 0 1
Fxc839_838 x839 0 Vx838 -416.31149371856
Cx839 x839 xm839 1.6602740464064e-14
Vx839 xm839 0 0
Gx839_2 x839 0 u2 0 3.47226538164996e-05
Rx840 x840 0 1
Fxc840_841 x840 0 Vx841 90.4352612427209
Cx840 x840 xm840 1.17924667928284e-12
Vx840 xm840 0 0
Gx840_2 x840 0 u2 0 -0.583193832252332
Rx841 x841 0 1
Fxc841_840 x841 0 Vx840 -2.57903242761661
Cx841 x841 xm841 1.17924667928284e-12
Vx841 xm841 0 0
Gx841_2 x841 0 u2 0 1.50407580496477
Rx842 x842 0 1
Fxc842_843 x842 0 Vx843 76.6151058397262
Cx842 x842 xm842 2.25551329603533e-13
Vx842 xm842 0 0
Gx842_2 x842 0 u2 0 -0.000961935158741434
Rx843 x843 0 1
Fxc843_842 x843 0 Vx842 -72.5569884446346
Cx843 x843 xm843 2.25551329603533e-13
Vx843 xm843 0 0
Gx843_2 x843 0 u2 0 0.06979511819729
Rx844 x844 0 1
Fxc844_845 x844 0 Vx845 1921.77776788372
Cx844 x844 xm844 3.84602500012975e-15
Vx844 xm844 0 0
Gx844_2 x844 0 u2 0 -1.80990219457151e-09
Rx845 x845 0 1
Fxc845_844 x845 0 Vx844 -9803.97529298039
Cx845 x845 xm845 3.84602500012975e-15
Vx845 xm845 0 0
Gx845_2 x845 0 u2 0 1.77442363982901e-05
Rx846 x846 0 1
Fxc846_847 x846 0 Vx847 15219.5253291423
Cx846 x846 xm846 9.27706506013979e-15
Vx846 xm846 0 0
Gx846_2 x846 0 u2 0 -2.46382987149046e-08
Rx847 x847 0 1
Fxc847_846 x847 0 Vx846 -214.696109142721
Cx847 x847 xm847 9.27706506013979e-15
Vx847 xm847 0 0
Gx847_2 x847 0 u2 0 5.28974686998613e-06
Rx848 x848 0 1
Fxc848_849 x848 0 Vx849 3400.29544354516
Cx848 x848 xm848 2.25851726135813e-15
Vx848 xm848 0 0
Gx848_2 x848 0 u2 0 -1.36437796648241e-09
Rx849 x849 0 1
Fxc849_848 x849 0 Vx848 -16342.0516313613
Cx849 x849 xm849 2.25851726135813e-15
Vx849 xm849 0 0
Gx849_2 x849 0 u2 0 2.22967351729472e-05
Rx850 x850 0 1
Fxc850_851 x850 0 Vx851 2117.34140011067
Cx850 x850 xm850 3.37035623112366e-15
Vx850 xm850 0 0
Gx850_2 x850 0 u2 0 -2.73280714065575e-09
Rx851 x851 0 1
Fxc851_850 x851 0 Vx850 -11895.9778828873
Cx851 x851 xm851 3.37035623112366e-15
Vx851 xm851 0 0
Gx851_2 x851 0 u2 0 3.25094133034371e-05
Rx852 x852 0 1
Fxc852_853 x852 0 Vx853 127.869920277283
Cx852 x852 xm852 1.88174133254326e-14
Vx852 xm852 0 0
Gx852_2 x852 0 u2 0 -2.20894852091485e-08
Rx853 x853 0 1
Fxc853_852 x853 0 Vx852 -6343.36616265804
Cx853 x853 xm853 1.88174133254326e-14
Vx853 xm853 0 0
Gx853_2 x853 0 u2 0 0.000140121693026248
Rx854 x854 0 1
Fxc854_855 x854 0 Vx855 1755.45429753074
Cx854 x854 xm854 1.207285936914e-14
Vx854 xm854 0 0
Gx854_2 x854 0 u2 0 -3.76911501062557e-08
Rx855 x855 0 1
Fxc855_854 x855 0 Vx854 -1130.40268606794
Cx855 x855 xm855 1.207285936914e-14
Vx855 xm855 0 0
Gx855_2 x855 0 u2 0 4.26061773211012e-05
Rx856 x856 0 1
Fxc856_857 x856 0 Vx857 4507.92221016949
Cx856 x856 xm856 1.59455172364102e-14
Vx856 xm856 0 0
Gx856_2 x856 0 u2 0 -4.29302862228671e-07
Rx857 x857 0 1
Fxc857_856 x857 0 Vx856 -254.590290772689
Cx857 x857 xm857 1.59455172364102e-14
Vx857 xm857 0 0
Gx857_2 x857 0 u2 0 0.000109296340524345
Rx858 x858 0 1
Fxc858_859 x858 0 Vx859 1547.44816345076
Cx858 x858 xm858 1.4256037936421e-14
Vx858 xm858 0 0
Gx858_2 x858 0 u2 0 -2.55970265627525e-07
Rx859 x859 0 1
Fxc859_858 x859 0 Vx858 -927.40393536027
Cx859 x859 xm859 1.4256037936421e-14
Vx859 xm859 0 0
Gx859_2 x859 0 u2 0 0.00023738783167818
Rx860 x860 0 1
Fxc860_861 x860 0 Vx861 57.0590012171719
Cx860 x860 xm860 1.54588556473979e-13
Vx860 xm860 0 0
Gx860_2 x860 0 u2 0 -4.1224508640184e-05
Rx861 x861 0 1
Fxc861_860 x861 0 Vx860 -217.748378182718
Cx861 x861 xm861 1.54588556473979e-13
Vx861 xm861 0 0
Gx861_2 x861 0 u2 0 0.0089765698977795
Rx862 x862 0 1
Fxc862_863 x862 0 Vx863 24723.718375191
Cx862 x862 xm862 1.36270438718843e-15
Vx862 xm862 0 0
Gx862_2 x862 0 u2 0 -2.96105151012464e-10
Rx863 x863 0 1
Fxc863_862 x863 0 Vx862 -6429.54979235673
Cx863 x863 xm863 1.36270438718843e-15
Vx863 xm863 0 0
Gx863_2 x863 0 u2 0 1.90382281220795e-06
Rx864 x864 0 1
Fxc864_865 x864 0 Vx865 222.008459848057
Cx864 x864 xm864 1.8842536609155e-14
Vx864 xm864 0 0
Gx864_2 x864 0 u2 0 -3.12935918377009e-08
Rx865 x865 0 1
Fxc865_864 x865 0 Vx864 -3762.01884295598
Cx865 x865 xm865 1.8842536609155e-14
Vx865 xm865 0 0
Gx865_2 x865 0 u2 0 0.000117727082157204
Rx866 x866 0 1
Fxc866_867 x866 0 Vx867 176.264808386761
Cx866 x866 xm866 2.58532363902921e-14
Vx866 xm866 0 0
Gx866_2 x866 0 u2 0 -8.22115047258298e-08
Rx867 x867 0 1
Fxc867_866 x867 0 Vx866 -2529.70492232687
Cx867 x867 xm867 2.58532363902921e-14
Vx867 xm867 0 0
Gx867_2 x867 0 u2 0 0.000207970848176831
Rx868 x868 0 1
Fxc868_869 x868 0 Vx869 8170.77518419377
Cx868 x868 xm868 4.40227995829476e-15
Vx868 xm868 0 0
Gx868_2 x868 0 u2 0 -2.91661001186959e-09
Rx869 x869 0 1
Fxc869_868 x869 0 Vx868 -1894.1525902487
Cx869 x869 xm869 4.40227995829476e-15
Vx869 xm869 0 0
Gx869_2 x869 0 u2 0 5.52450440872808e-06
Rx870 x870 0 1
Fxc870_871 x870 0 Vx871 603.170742581347
Cx870 x870 xm870 2.0912663085398e-14
Vx870 xm870 0 0
Gx870_2 x870 0 u2 0 -8.4346709754617e-08
Rx871 x871 0 1
Fxc871_870 x871 0 Vx870 -1146.35910168148
Cx871 x871 xm871 2.0912663085398e-14
Vx871 xm871 0 0
Gx871_2 x871 0 u2 0 9.66916184240915e-05
Rx872 x872 0 1
Fxc872_873 x872 0 Vx873 730.070519195499
Cx872 x872 xm872 6.45713973054353e-15
Vx872 xm872 0 0
Gx872_2 x872 0 u2 0 -2.44990689398813e-09
Rx873 x873 0 1
Fxc873_872 x873 0 Vx872 -10017.1516461714
Cx873 x873 xm873 6.45713973054353e-15
Vx873 xm873 0 0
Gx873_2 x873 0 u2 0 2.454108887608e-05
Rx874 x874 0 1
Fxc874_875 x874 0 Vx875 5182.56835629346
Cx874 x874 xm874 7.88540425403586e-15
Vx874 xm874 0 0
Gx874_2 x874 0 u2 0 -1.01152303736804e-08
Rx875 x875 0 1
Fxc875_874 x875 0 Vx874 -951.571775973863
Cx875 x875 xm875 7.88540425403586e-15
Vx875 xm875 0 0
Gx875_2 x875 0 u2 0 9.62536773106778e-06
Rx876 x876 0 1
Fxc876_877 x876 0 Vx877 46.5148157503785
Cx876 x876 xm876 1.62084283086177e-13
Vx876 xm876 0 0
Gx876_2 x876 0 u2 0 -2.37858331327793e-05
Rx877 x877 0 1
Fxc877_876 x877 0 Vx876 -267.354608863644
Cx877 x877 xm877 1.62084283086177e-13
Vx877 xm877 0 0
Gx877_2 x877 0 u2 0 0.00635925211371011
Rx878 x878 0 1
Fxc878_879 x878 0 Vx879 813.940595162096
Cx878 x878 xm878 5.31549963067726e-14
Vx878 xm878 0 0
Gx878_2 x878 0 u2 0 -1.597258678323e-06
Rx879 x879 0 1
Fxc879_878 x879 0 Vx878 -135.097678885803
Cx879 x879 xm879 5.31549963067726e-14
Vx879 xm879 0 0
Gx879_2 x879 0 u2 0 0.000215785940021642
Rx880 x880 0 1
Fxc880_881 x880 0 Vx881 377.959888195475
Cx880 x880 xm880 1.78816112180161e-14
Vx880 xm880 0 0
Gx880_2 x880 0 u2 0 -3.54231905087853e-08
Rx881 x881 0 1
Fxc881_880 x881 0 Vx880 -2560.56460017476
Cx881 x881 xm881 1.78816112180161e-14
Vx881 xm881 0 0
Gx881_2 x881 0 u2 0 9.07033676420419e-05
Rx882 x882 0 1
Fxc882_883 x882 0 Vx883 1885.27822840143
Cx882 x882 xm882 7.76754927887759e-15
Vx882 xm882 0 0
Gx882_2 x882 0 u2 0 -5.53905769111327e-09
Rx883 x883 0 1
Fxc883_882 x883 0 Vx882 -2747.28042669389
Cx883 x883 xm883 7.7675492788776e-15
Vx883 xm883 0 0
Gx883_2 x883 0 u2 0 1.52173447771237e-05
Rx884 x884 0 1
Fxc884_885 x884 0 Vx885 48529.8782933035
Cx884 x884 xm884 1.25557410678191e-15
Vx884 xm884 0 0
Gx884_2 x884 0 u2 0 -5.87433275684117e-11
Rx885 x885 0 1
Fxc885_884 x885 0 Vx884 -4109.7287529175
Cx885 x885 xm885 1.25557410678191e-15
Vx885 xm885 0 0
Gx885_2 x885 0 u2 0 2.41419142349953e-07
Rx886 x886 0 1
Fxc886_887 x886 0 Vx887 482.378013054463
Cx886 x886 xm886 1.63787697489454e-14
Vx886 xm886 0 0
Gx886_2 x886 0 u2 0 -2.45576214512506e-08
Rx887 x887 0 1
Fxc887_886 x887 0 Vx886 -2527.67699045898
Cx887 x887 xm887 1.63787697489454e-14
Vx887 xm887 0 0
Gx887_2 x887 0 u2 0 6.20737346827279e-05
Rx888 x888 0 1
Fxc888_889 x888 0 Vx889 3404.69443339039
Cx888 x888 xm888 1.19981261746115e-15
Vx888 xm888 0 0
Gx888_2 x888 0 u2 0 -3.86890396666103e-11
Rx889 x889 0 1
Fxc889_888 x889 0 Vx888 -64529.8857673097
Cx889 x889 xm889 1.19981261746115e-15
Vx889 xm889 0 0
Gx889_2 x889 0 u2 0 2.49659931013328e-06
Rx890 x890 0 1
Fxc890_891 x890 0 Vx891 33003.1514471578
Cx890 x890 xm890 6.90011418477151e-16
Vx890 xm890 0 0
Gx890_2 x890 0 u2 0 -7.6120518018319e-10
Rx891 x891 0 1
Fxc891_890 x891 0 Vx890 -20721.6257270503
Cx891 x891 xm891 6.90011418477151e-16
Vx891 xm891 0 0
Gx891_2 x891 0 u2 0 1.57734088452479e-05
Rx892 x892 0 1
Fxc892_893 x892 0 Vx893 54395.6929100173
Cx892 x892 xm892 1.91401504019507e-14
Vx892 xm892 0 0
Gx892_2 x892 0 u2 0 -1.1143950123431e-07
Rx893 x893 0 1
Fxc893_892 x893 0 Vx892 -16.1640053968643
Cx893 x893 xm893 1.91401504019507e-14
Vx893 xm893 0 0
Gx893_2 x893 0 u2 0 1.80130869937525e-06
Rx894 x894 0 1
Fxc894_895 x894 0 Vx895 442.226084175693
Cx894 x894 xm894 2.78471100161717e-14
Vx894 xm894 0 0
Gx894_2 x894 0 u2 0 -1.86024354967913e-07
Rx895 x895 0 1
Fxc895_894 x895 0 Vx894 -942.881099206962
Cx895 x895 xm895 2.78471100161717e-14
Vx895 xm895 0 0
Gx895_2 x895 0 u2 0 0.000175398848291411
Rx896 x896 0 1
Fxc896_897 x896 0 Vx897 5220.03110549995
Cx896 x896 xm896 7.87159377020613e-15
Vx896 xm896 0 0
Gx896_2 x896 0 u2 0 -9.67405371781818e-09
Rx897 x897 0 1
Fxc897_896 x897 0 Vx896 -984.959492791397
Cx897 x897 xm897 7.87159377020614e-15
Vx897 xm897 0 0
Gx897_2 x897 0 u2 0 9.52855104313892e-06
Rx898 x898 0 1
Fxc898_899 x898 0 Vx899 5.618557622684
Cx898 x898 xm898 1.06813886291274e-12
Vx898 xm898 0 0
Gx898_2 x898 0 u2 0 -0.087019371453461
Rx899 x899 0 1
Fxc899_898 x899 0 Vx898 -52.7418861736944
Cx899 x899 xm899 1.06813886291274e-12
Vx899 xm899 0 0
Gx899_2 x899 0 u2 0 4.58956578410488
Rx900 x900 0 1
Fxc900_901 x900 0 Vx901 76584.8940565089
Cx900 x900 xm900 5.25955260177112e-15
Vx900 xm900 0 0
Gx900_2 x900 0 u2 0 -2.88830282124005e-09
Rx901 x901 0 1
Fxc901_900 x901 0 Vx900 -155.313739876454
Cx901 x901 xm901 5.25955260177112e-15
Vx901 xm901 0 0
Gx901_2 x901 0 u2 0 4.48593113062507e-07
Rx902 x902 0 1
Fxc902_903 x902 0 Vx903 441.872182266179
Cx902 x902 xm902 2.76085682247672e-14
Vx902 xm902 0 0
Gx902_2 x902 0 u2 0 -1.32088490162406e-07
Rx903 x903 0 1
Fxc903_902 x903 0 Vx902 -984.596532880146
Cx903 x903 xm903 2.76085682247672e-14
Vx903 xm903 0 0
Gx903_2 x903 0 u2 0 0.000130053869447279
Rx904 x904 0 1
Fxc904_905 x904 0 Vx905 234.113892659305
Cx904 x904 xm904 1.46519190092729e-14
Vx904 xm904 0 0
Gx904_2 x904 0 u2 0 -8.84754912612056e-09
Rx905 x905 0 1
Fxc905_904 x905 0 Vx904 -6640.82702000552
Cx905 x905 xm905 1.46519190092729e-14
Vx905 xm905 0 0
Gx905_2 x905 0 u2 0 5.87550432975676e-05
Rx906 x906 0 1
Fxc906_907 x906 0 Vx907 2239.06515216328
Cx906 x906 xm906 2.19788949285279e-14
Vx906 xm906 0 0
Gx906_2 x906 0 u2 0 -1.08111289494745e-07
Rx907 x907 0 1
Fxc907_906 x907 0 Vx906 -311.183105419374
Cx907 x907 xm907 2.19788949285279e-14
Vx907 xm907 0 0
Gx907_2 x907 0 u2 0 3.36424067958678e-05
Rx908 x908 0 1
Fxc908_909 x908 0 Vx909 750.114431051507
Cx908 x908 xm908 8.20375533487514e-14
Vx908 xm908 0 0
Gx908_2 x908 0 u2 0 -4.27619568501889e-06
Rx909 x909 0 1
Fxc909_908 x909 0 Vx908 -67.3355989831271
Cx909 x909 xm909 8.20375533487514e-14
Vx909 xm909 0 0
Gx909_2 x909 0 u2 0 0.000287940197819811
Rx910 x910 0 1
Fxc910_911 x910 0 Vx911 2532.37423032255
Cx910 x910 xm910 7.51272397073094e-15
Vx910 xm910 0 0
Gx910_2 x910 0 u2 0 -5.82110520200593e-09
Rx911 x911 0 1
Fxc911_910 x911 0 Vx910 -2384.62854254448
Cx911 x911 xm911 7.51272397073094e-15
Vx911 xm911 0 0
Gx911_2 x911 0 u2 0 1.38811736138575e-05
Rx912 x912 0 1
Fxc912_913 x912 0 Vx913 985.222260913355
Cx912 x912 xm912 1.25924088295157e-14
Vx912 xm912 0 0
Gx912_2 x912 0 u2 0 -1.63704363292285e-08
Rx913 x913 0 1
Fxc913_912 x913 0 Vx912 -2360.74888854806
Cx913 x913 xm913 1.25924088295157e-14
Vx913 xm913 0 0
Gx913_2 x913 0 u2 0 3.8646489369273e-05
Rx914 x914 0 1
Fxc914_915 x914 0 Vx915 353.441075041497
Cx914 x914 xm914 3.99671423619986e-14
Vx914 xm914 0 0
Gx914_2 x914 0 u2 0 -3.44836075634036e-07
Rx915 x915 0 1
Fxc915_914 x915 0 Vx914 -649.571514967075
Cx915 x915 xm915 3.99671423619986e-14
Vx915 xm915 0 0
Gx915_2 x915 0 u2 0 0.000223995692064902
Rx916 x916 0 1
Fxc916_917 x916 0 Vx917 1822.21575339883
Cx916 x916 xm916 4.75295253243805e-15
Vx916 xm916 0 0
Gx916_2 x916 0 u2 0 -2.63577542158311e-09
Rx917 x917 0 1
Fxc917_916 x917 0 Vx916 -8381.46521596228
Cx917 x917 xm917 4.75295253243805e-15
Vx917 xm917 0 0
Gx917_2 x917 0 u2 0 2.20916600130872e-05
Rx918 x918 0 1
Fxc918_919 x918 0 Vx919 371.787347184655
Cx918 x918 xm918 3.41070990725561e-14
Vx918 xm918 0 0
Gx918_2 x918 0 u2 0 -1.84049381307143e-07
Rx919 x919 0 1
Fxc919_918 x919 0 Vx918 -801.787616879464
Cx919 x919 xm919 3.41070990725561e-14
Vx919 xm919 0 0
Gx919_2 x919 0 u2 0 0.000147568514826394
Rx920 x920 0 1
Fxc920_921 x920 0 Vx921 2174.81451507683
Cx920 x920 xm920 9.91623794270551e-15
Vx920 xm920 0 0
Gx920_2 x920 0 u2 0 -1.29932499865672e-08
Rx921 x921 0 1
Fxc921_920 x921 0 Vx920 -1631.34741653125
Cx921 x921 xm921 9.91623794270551e-15
Vx921 xm921 0 0
Gx921_2 x921 0 u2 0 2.11965047979312e-05
Rx922 x922 0 1
Fxc922_923 x922 0 Vx923 209.439421905225
Cx922 x922 xm922 2.22232201775079e-14
Vx922 xm922 0 0
Gx922_2 x922 0 u2 0 -2.92115832519093e-08
Rx923 x923 0 1
Fxc923_922 x923 0 Vx922 -3512.03650866934
Cx923 x923 xm923 2.22232201775079e-14
Vx923 xm923 0 0
Gx923_2 x923 0 u2 0 0.000102592146856739
Rx924 x924 0 1
Fxc924_925 x924 0 Vx925 4432.48862054229
Cx924 x924 xm924 5.17797017606527e-15
Vx924 xm924 0 0
Gx924_2 x924 0 u2 0 -2.16337717018969e-09
Rx925 x925 0 1
Fxc925_924 x925 0 Vx924 -2957.63385008778
Cx925 x925 xm925 5.17797017606527e-15
Vx925 xm925 0 0
Gx925_2 x925 0 u2 0 6.39847754906015e-06
Rx926 x926 0 1
Fxc926_927 x926 0 Vx927 198.06283356188
Cx926 x926 xm926 4.46596707298567e-14
Vx926 xm926 0 0
Gx926_2 x926 0 u2 0 -4.16398122175432e-07
Rx927 x927 0 1
Fxc927_926 x927 0 Vx926 -902.555971169995
Cx927 x927 xm927 4.46596707298567e-14
Vx927 xm927 0 0
Gx927_2 x927 0 u2 0 0.000375822611553409
Rx928 x928 0 1
Fxc928_929 x928 0 Vx929 394.775883842956
Cx928 x928 xm928 1.25147099405371e-14
Vx928 xm928 0 0
Gx928_2 x928 0 u2 0 -7.93652929105126e-09
Rx929 x929 0 1
Fxc929_928 x929 0 Vx928 -5846.15772382472
Cx929 x929 xm929 1.25147099405371e-14
Vx929 xm929 0 0
Gx929_2 x929 0 u2 0 4.63982020152405e-05
Rx930 x930 0 1
Fxc930_931 x930 0 Vx931 27968.4767076373
Cx930 x930 xm930 3.07868023406084e-14
Vx930 xm930 0 0
Gx930_2 x930 0 u2 0 -3.61694566677464e-07
Rx931 x931 0 1
Fxc931_930 x931 0 Vx930 -13.5278441690684
Cx931 x931 xm931 3.07868023406084e-14
Vx931 xm931 0 0
Gx931_2 x931 0 u2 0 4.89294773481144e-06
Rx932 x932 0 1
Fxc932_933 x932 0 Vx933 1366.07700198898
Cx932 x932 xm932 5.4585280782342e-15
Vx932 xm932 0 0
Gx932_2 x932 0 u2 0 -1.71077207485317e-09
Rx933 x933 0 1
Fxc933_932 x933 0 Vx932 -8763.1913119305
Cx933 x933 xm933 5.4585280782342e-15
Vx933 xm933 0 0
Gx933_2 x933 0 u2 0 1.49918229830466e-05
Rx934 x934 0 1
Fxc934_935 x934 0 Vx935 18.0353919338892
Cx934 x934 xm934 2.51329289587019e-12
Vx934 xm934 0 0
Gx934_2 x934 0 u2 0 -3.79660896437117
Rx935 x935 0 1
Fxc935_934 x935 0 Vx934 -3.75811865469954
Cx935 x935 xm935 2.51329289587019e-12
Vx935 xm935 0 0
Gx935_2 x935 0 u2 0 14.2681069736028
Rx936 x936 0 1
Fxc936_937 x936 0 Vx937 80.6224231967355
Cx936 x936 xm936 3.57049647256315e-13
Vx936 xm936 0 0
Gx936_2 x936 0 u2 0 -0.000506515516249674
Rx937 x937 0 1
Fxc937_936 x937 0 Vx936 -39.9726183030067
Cx937 x937 xm937 3.57049647256315e-13
Vx937 xm937 0 0
Gx937_2 x937 0 u2 0 0.0202467513955986
Rx938 x938 0 1
Fxc938_939 x938 0 Vx939 603.4590823449
Cx938 x938 xm938 4.5035441503013e-14
Vx938 xm938 0 0
Gx938_2 x938 0 u2 0 -5.97666498618081e-07
Rx939 x939 0 1
Fxc939_938 x939 0 Vx938 -303.351510767652
Cx939 x939 xm939 4.5035441503013e-14
Vx939 xm939 0 0
Gx939_2 x939 0 u2 0 0.000181303035291008
Rx940 x940 0 1
Fxc940_941 x940 0 Vx941 1727.33129617615
Cx940 x940 xm940 8.56467633357547e-15
Vx940 xm940 0 0
Gx940_2 x940 0 u2 0 -8.81640431328412e-09
Rx941 x941 0 1
Fxc941_940 x941 0 Vx940 -2958.44455508609
Cx941 x941 xm941 8.56467633357547e-15
Vx941 xm941 0 0
Gx941_2 x941 0 u2 0 2.6082843336073e-05
Rx942 x942 0 1
Fxc942_943 x942 0 Vx943 90.7659929353874
Cx942 x942 xm942 8.27372304605411e-14
Vx942 xm942 0 0
Gx942_2 x942 0 u2 0 -8.47690579013902e-07
Rx943 x943 0 1
Fxc943_942 x943 0 Vx942 -648.325093622117
Cx943 x943 xm943 8.27372304605411e-14
Vx943 xm943 0 0
Gx943_2 x943 0 u2 0 0.000549579074001775
Rx944 x944 0 1
Fxc944_945 x944 0 Vx945 1086.92406503906
Cx944 x944 xm944 1.66721817308413e-14
Vx944 xm944 0 0
Gx944_2 x944 0 u2 0 -3.9337783595517e-08
Rx945 x945 0 1
Fxc945_944 x945 0 Vx944 -1247.25734073378
Cx945 x945 xm945 1.66721817308413e-14
Vx945 xm945 0 0
Gx945_2 x945 0 u2 0 4.90643393577055e-05
Rx946 x946 0 1
Fxc946_947 x946 0 Vx947 1574.62365002861
Cx946 x946 xm946 7.0052963467164e-14
Vx946 xm946 0 0
Gx946_2 x946 0 u2 0 -3.1333811152908e-06
Rx947 x947 0 1
Fxc947_946 x947 0 Vx946 -48.8622549359032
Cx947 x947 xm947 7.00529634671639e-14
Vx947 xm947 0 0
Gx947_2 x947 0 u2 0 0.000153104066866684
Rx948 x948 0 1
Fxc948_949 x948 0 Vx949 842804.932016304
Cx948 x948 xm948 1.10677227211622e-16
Vx948 xm948 0 0
Gx948_2 x948 0 u2 0 -1.27907379888214e-11
Rx949 x949 0 1
Fxc949_948 x949 0 Vx948 -38909.7733336474
Cx949 x949 xm949 1.10677227211622e-16
Vx949 xm949 0 0
Gx949_2 x949 0 u2 0 4.97684715915113e-07
Rx950 x950 0 1
Fxc950_951 x950 0 Vx951 8926.99017004506
Cx950 x950 xm950 1.5846769699005e-14
Vx950 xm950 0 0
Gx950_2 x950 0 u2 0 -2.68295365849138e-08
Rx951 x951 0 1
Fxc951_950 x951 0 Vx950 -177.292051713135
Cx951 x951 xm951 1.5846769699005e-14
Vx951 xm951 0 0
Gx951_2 x951 0 u2 0 4.75666358765198e-06
Rx952 x952 0 1
Fxc952_953 x952 0 Vx953 890.244484805097
Cx952 x952 xm952 4.12031373830175e-14
Vx952 xm952 0 0
Gx952_2 x952 0 u2 0 -1.0630555057862e-06
Rx953 x953 0 1
Fxc953_952 x953 0 Vx952 -254.81230161624
Cx953 x953 xm953 4.12031373830175e-14
Vx953 xm953 0 0
Gx953_2 x953 0 u2 0 0.000270879620175196
Rx954 x954 0 1
Fxc954_955 x954 0 Vx955 1731.91381828514
Cx954 x954 xm954 1.43266280058829e-14
Vx954 xm954 0 0
Gx954_2 x954 0 u2 0 -2.74603684506172e-08
Rx955 x955 0 1
Fxc955_954 x955 0 Vx954 -1077.20255022272
Cx955 x955 xm955 1.43266280058829e-14
Vx955 xm955 0 0
Gx955_2 x955 0 u2 0 2.95803789250604e-05
Rx956 x956 0 1
Fxc956_957 x956 0 Vx957 294.98398496282
Cx956 x956 xm956 9.37589835741656e-14
Vx956 xm956 0 0
Gx956_2 x956 0 u2 0 -8.2787723349726e-06
Rx957 x957 0 1
Fxc957_956 x957 0 Vx956 -149.602993024203
Cx957 x957 xm957 9.37589835741656e-14
Vx957 xm957 0 0
Gx957_2 x957 0 u2 0 0.00123852911987787
Rx958 x958 0 1
Fxc958_959 x958 0 Vx959 2146.01426892351
Cx958 x958 xm958 2.94431934184726e-15
Vx958 xm958 0 0
Gx958_2 x958 0 u2 0 -1.23330684204259e-10
Rx959 x959 0 1
Fxc959_958 x959 0 Vx958 -20990.5196704473
Cx959 x959 xm959 2.94431934184726e-15
Vx959 xm959 0 0
Gx959_2 x959 0 u2 0 2.58877515275922e-06
Rx960 x960 0 1
Fxc960_961 x960 0 Vx961 127606.83195335
Cx960 x960 xm960 1.38008738267159e-16
Vx960 xm960 0 0
Gx960_2 x960 0 u2 0 -6.92416359582259e-11
Rx961 x961 0 1
Fxc961_960 x961 0 Vx960 -162101.840431999
Cx961 x961 xm961 1.38008738267159e-16
Vx961 xm961 0 0
Gx961_2 x961 0 u2 0 1.12241966233509e-05
Rx962 x962 0 1
Fxc962_963 x962 0 Vx963 184.422161853856
Cx962 x962 xm962 3.31616743972311e-14
Vx962 xm962 0 0
Gx962_2 x962 0 u2 0 -1.92067186572256e-07
Rx963 x963 0 1
Fxc963_962 x963 0 Vx962 -1906.69005516502
Cx963 x963 xm963 3.31616743972311e-14
Vx963 xm963 0 0
Gx963_2 x963 0 u2 0 0.000366212594560846
Rx964 x964 0 1
Fxc964_965 x964 0 Vx965 22.3433589997169
Cx964 x964 xm964 6.8171023360865e-13
Vx964 xm964 0 0
Gx964_2 x964 0 u2 0 -0.0114551334864184
Rx965 x965 0 1
Fxc965_964 x965 0 Vx964 -41.6969609809194
Cx965 x965 xm965 6.8171023360865e-13
Vx965 xm965 0 0
Gx965_2 x965 0 u2 0 0.47764425401441
Rx966 x966 0 1
Fxc966_967 x966 0 Vx967 9353.88063386068
Cx966 x966 xm966 1.6412792293327e-15
Vx966 xm966 0 0
Gx966_2 x966 0 u2 0 -4.64247929762518e-10
Rx967 x967 0 1
Fxc967_966 x967 0 Vx966 -16130.415652273
Cx967 x967 xm967 1.6412792293327e-15
Vx967 xm967 0 0
Gx967_2 x967 0 u2 0 7.48851207277666e-06
Rx968 x968 0 1
Fxc968_969 x968 0 Vx969 97.7741336245745
Cx968 x968 xm968 2.0277279276718e-14
Vx968 xm968 0 0
Gx968_2 x968 0 u2 0 -5.84229909621269e-09
Rx969 x969 0 1
Fxc969_968 x969 0 Vx968 -10860.3239755057
Cx969 x969 xm969 2.0277279276718e-14
Vx969 xm969 0 0
Gx969_2 x969 0 u2 0 6.3449260946674e-05
Rx970 x970 0 1
Fxc970_971 x970 0 Vx971 1877.20718852291
Cx970 x970 xm970 9.54778893264496e-15
Vx970 xm970 0 0
Gx970_2 x970 0 u2 0 -6.83633260292491e-09
Rx971 x971 0 1
Fxc971_970 x971 0 Vx970 -2386.81092912641
Cx971 x971 xm971 9.54778893264496e-15
Vx971 xm971 0 0
Gx971_2 x971 0 u2 0 1.63170333718043e-05
Rx972 x972 0 1
Fxc972_973 x972 0 Vx973 1032.75941035992
Cx972 x972 xm972 1.33797401275805e-14
Vx972 xm972 0 0
Gx972_2 x972 0 u2 0 -8.46410005713732e-09
Rx973 x973 0 1
Fxc973_972 x973 0 Vx972 -2229.80625568951
Cx973 x973 xm973 1.33797401275805e-14
Vx973 xm973 0 0
Gx973_2 x973 0 u2 0 1.88733032561867e-05
Rx974 x974 0 1
Fxc974_975 x974 0 Vx975 41399.0565697948
Cx974 x974 xm974 8.17600979330828e-15
Vx974 xm974 0 0
Gx974_2 x974 0 u2 0 -6.95045437437488e-09
Rx975 x975 0 1
Fxc975_974 x975 0 Vx974 -151.256126978571
Cx975 x975 xm975 8.17600979330828e-15
Vx975 xm975 0 0
Gx975_2 x975 0 u2 0 1.05129880940921e-06
Rx976 x976 0 1
Fxc976_977 x976 0 Vx977 887.076179277472
Cx976 x976 xm976 1.96425850879399e-14
Vx976 xm976 0 0
Gx976_2 x976 0 u2 0 -3.19050537955219e-08
Rx977 x977 0 1
Fxc977_976 x977 0 Vx976 -1259.66151506927
Cx977 x977 xm977 1.96425850879399e-14
Vx977 xm977 0 0
Gx977_2 x977 0 u2 0 4.01895684024338e-05
Rx978 x978 0 1
Fxc978_979 x978 0 Vx979 904.387819043909
Cx978 x978 xm978 1.88286053329382e-14
Vx978 xm978 0 0
Gx978_2 x978 0 u2 0 -3.54463653109283e-08
Rx979 x979 0 1
Fxc979_978 x979 0 Vx978 -1356.38135680894
Cx979 x979 xm979 1.88286053329382e-14
Vx979 xm979 0 0
Gx979_2 x979 0 u2 0 4.80787890743823e-05
Rx980 x980 0 1
Fxc980_981 x980 0 Vx981 3216.74965143391
Cx980 x980 xm980 1.88018559993273e-14
Vx980 xm980 0 0
Gx980_2 x980 0 u2 0 -5.02541620380387e-08
Rx981 x981 0 1
Fxc981_980 x981 0 Vx980 -376.051609572161
Cx981 x981 xm981 1.88018559993273e-14
Vx981 xm981 0 0
Gx981_2 x981 0 u2 0 1.88981585221046e-05
Rx982 x982 0 1
Fxc982_983 x982 0 Vx983 5740.76490231102
Cx982 x982 xm982 1.24637336182944e-15
Vx982 xm982 0 0
Gx982_2 x982 0 u2 0 -2.54784723603567e-10
Rx983 x983 0 1
Fxc983_982 x983 0 Vx982 -46696.7867368399
Cx983 x983 xm983 1.24637336182943e-15
Vx983 xm983 0 0
Gx983_2 x983 0 u2 0 1.18976279019205e-05
Rx984 x984 0 1
Fxc984_985 x984 0 Vx985 2223.31233356045
Cx984 x984 xm984 9.701039005748e-15
Vx984 xm984 0 0
Gx984_2 x984 0 u2 0 -1.12886514955727e-08
Rx985 x985 0 1
Fxc985_984 x985 0 Vx984 -2017.47802443671
Cx985 x985 xm985 9.701039005748e-15
Vx985 xm985 0 0
Gx985_2 x985 0 u2 0 2.27746063178426e-05
Rx986 x986 0 1
Fxc986_987 x986 0 Vx987 750.492731303233
Cx986 x986 xm986 2.77515669599418e-14
Vx986 xm986 0 0
Gx986_2 x986 0 u2 0 -1.00572744627923e-07
Rx987 x987 0 1
Fxc987_986 x987 0 Vx986 -734.573437844736
Cx987 x987 xm987 2.77515669599418e-14
Vx987 xm987 0 0
Gx987_2 x987 0 u2 0 7.3878066774814e-05
Rx988 x988 0 1
Fxc988_989 x988 0 Vx989 31.5120562158234
Cx988 x988 xm988 1.90385021922328e-12
Vx988 xm988 0 0
Gx988_2 x988 0 u2 0 -1.05787127404968
Rx989 x989 0 1
Fxc989_988 x989 0 Vx988 -4.15315854255383
Cx989 x989 xm989 1.90385021922328e-12
Vx989 xm989 0 0
Gx989_2 x989 0 u2 0 4.39350711874173
Rx990 x990 0 1
Fxc990_991 x990 0 Vx991 126.123865782952
Cx990 x990 xm990 4.13080608699608e-13
Vx990 xm990 0 0
Gx990_2 x990 0 u2 0 -0.00290100913361198
Rx991 x991 0 1
Fxc991_990 x991 0 Vx990 -21.8738925891598
Cx991 x991 xm991 4.13080608699608e-13
Vx991 xm991 0 0
Gx991_2 x991 0 u2 0 0.0634563621887998
Rx992 x992 0 1
Fxc992_993 x992 0 Vx993 7.4626585353331
Cx992 x992 xm992 3.88335929258945e-13
Vx992 xm992 0 0
Gx992_2 x992 0 u2 0 -0.000741651051826747
Rx993 x993 0 1
Fxc993_992 x993 0 Vx992 -407.387970315477
Cx993 x993 xm993 3.88335929258946e-13
Vx993 xm993 0 0
Gx993_2 x993 0 u2 0 0.302139716686037
Rx994 x994 0 1
Fxc994_995 x994 0 Vx995 93.3363626355421
Cx994 x994 xm994 2.37282917151686e-13
Vx994 xm994 0 0
Gx994_2 x994 0 u2 0 -0.000379824149638761
Rx995 x995 0 1
Fxc995_994 x995 0 Vx994 -86.6527515050668
Cx995 x995 xm995 2.37282917151686e-13
Vx995 xm995 0 0
Gx995_2 x995 0 u2 0 0.0329128076542709
Rx996 x996 0 1
Fxc996_997 x996 0 Vx997 605.482578464241
Cx996 x996 xm996 1.91607970073068e-14
Vx996 xm996 0 0
Gx996_2 x996 0 u2 0 -1.96448387782998e-08
Rx997 x997 0 1
Fxc997_996 x997 0 Vx996 -1995.2465005569
Cx997 x997 xm997 1.91607970073068e-14
Vx997 xm997 0 0
Gx997_2 x997 0 u2 0 3.91962958264072e-05
Rx998 x998 0 1
Fxc998_999 x998 0 Vx999 180159.028077109
Cx998 x998 xm998 2.33334731840831e-14
Vx998 xm998 0 0
Gx998_2 x998 0 u2 0 -9.17975584779295e-08
Rx999 x999 0 1
Fxc999_998 x999 0 Vx998 -4.76014404799589
Cx999 x999 xm999 2.33334731840831e-14
Vx999 xm999 0 0
Gx999_2 x999 0 u2 0 4.36969601609271e-07
Rx1000 x1000 0 1
Fxc1000_1001 x1000 0 Vx1001 8021.78672121851
Cx1000 x1000 xm1000 2.2448315996525e-14
Vx1000 xm1000 0 0
Gx1000_2 x1000 0 u2 0 -8.95343877380737e-08
Rx1001 x1001 0 1
Fxc1001_1000 x1001 0 Vx1000 -114.920717799488
Cx1001 x1001 xm1001 2.2448315996525e-14
Vx1001 xm1001 0 0
Gx1001_2 x1001 0 u2 0 1.02893561065971e-05
Rx1002 x1002 0 1
Fxc1002_1003 x1002 0 Vx1003 461.353255388419
Cx1002 x1002 xm1002 5.50128571655933e-15
Vx1002 xm1002 0 0
Gx1002_2 x1002 0 u2 0 -3.24435712963443e-10
Rx1003 x1003 0 1
Fxc1003_1002 x1003 0 Vx1002 -32995.3879375282
Cx1003 x1003 xm1003 5.50128571655933e-15
Vx1003 xm1003 0 0
Gx1003_2 x1003 0 u2 0 1.07048822100174e-05
Rx1004 x1004 0 1
Fxc1004_1005 x1004 0 Vx1005 556.011051948472
Cx1004 x1004 xm1004 5.82585824065102e-14
Vx1004 xm1004 0 0
Gx1004_2 x1004 0 u2 0 -1.07927473720351e-06
Rx1005 x1005 0 1
Fxc1005_1004 x1005 0 Vx1004 -239.935193423816
Cx1005 x1005 xm1005 5.82585824065102e-14
Vx1005 xm1005 0 0
Gx1005_2 x1005 0 u2 0 0.000258955992828361
Rx1006 x1006 0 1
Fxc1006_1007 x1006 0 Vx1007 2015.44261340264
Cx1006 x1006 xm1006 4.64126067377759e-16
Vx1006 xm1006 0 0
Gx1006_2 x1006 0 u2 0 -8.37459256821118e-12
Rx1007 x1007 0 1
Fxc1007_1006 x1007 0 Vx1006 -1040345.89123581
Cx1007 x1007 xm1007 4.64126067377759e-16
Vx1007 xm1007 0 0
Gx1007_2 x1007 0 u2 0 8.71247296911247e-06
Rx1008 x1008 0 1
Fxc1008_1009 x1008 0 Vx1009 9903.26927416426
Cx1008 x1008 xm1008 4.79316217773287e-15
Vx1008 xm1008 0 0
Gx1008_2 x1008 0 u2 0 -2.53204579493926e-09
Rx1009 x1009 0 1
Fxc1009_1008 x1009 0 Vx1008 -1964.02612600966
Cx1009 x1009 xm1009 4.79316217773287e-15
Vx1009 xm1009 0 0
Gx1009_2 x1009 0 u2 0 4.97300409351361e-06
Rx1010 x1010 0 1
Fxc1010_1011 x1010 0 Vx1011 2.16336345065091
Cx1010 x1010 xm1010 4.88202959865766e-12
Vx1010 xm1010 0 0
Gx1010_2 x1010 0 u2 0 -1.52574856885853
Rx1011 x1011 0 1
Fxc1011_1010 x1011 0 Vx1010 -11.259372503232
Cx1011 x1011 xm1011 4.88202959865766e-12
Vx1011 xm1011 0 0
Gx1011_2 x1011 0 u2 0 17.1789714830514
Rx1012 x1012 0 1
Fxc1012_1013 x1012 0 Vx1013 4435.24951021907
Cx1012 x1012 xm1012 3.10944035248846e-15
Vx1012 xm1012 0 0
Gx1012_2 x1012 0 u2 0 -3.08525946249681e-10
Rx1013 x1013 0 1
Fxc1013_1012 x1013 0 Vx1012 -11051.9646966392
Cx1013 x1013 xm1013 3.10944035248846e-15
Vx1013 xm1013 0 0
Gx1013_2 x1013 0 u2 0 3.40981786594868e-06
Rx1014 x1014 0 1
Fxc1014_1015 x1014 0 Vx1015 700.2631577964
Cx1014 x1014 xm1014 2.0409012950473e-14
Vx1014 xm1014 0 0
Gx1014_2 x1014 0 u2 0 -4.04560487950749e-08
Rx1015 x1015 0 1
Fxc1015_1014 x1015 0 Vx1014 -1641.7894920117
Cx1015 x1015 xm1015 2.0409012950473e-14
Vx1015 xm1015 0 0
Gx1015_2 x1015 0 u2 0 6.64203158000668e-05
Rx1016 x1016 0 1
Fxc1016_1017 x1016 0 Vx1017 1230.92615649877
Cx1016 x1016 xm1016 4.35243189785395e-14
Vx1016 xm1016 0 0
Gx1016_2 x1016 0 u2 0 -1.12618380598557e-06
Rx1017 x1017 0 1
Fxc1017_1016 x1017 0 Vx1016 -207.286626371561
Cx1017 x1017 xm1017 4.35243189785395e-14
Vx1017 xm1017 0 0
Gx1017_2 x1017 0 u2 0 0.000233442841817032
Rx1018 x1018 0 1
Fxc1018_1019 x1018 0 Vx1019 427.95043321454
Cx1018 x1018 xm1018 4.3066796599514e-14
Vx1018 xm1018 0 0
Gx1018_2 x1018 0 u2 0 -6.88611855476646e-07
Rx1019 x1019 0 1
Fxc1019_1018 x1019 0 Vx1018 -606.702127687178
Cx1019 x1019 xm1019 4.30667965995139e-14
Vx1019 xm1019 0 0
Gx1019_2 x1019 0 u2 0 0.000417782277868297
Rx1020 x1020 0 1
Fxc1020_1021 x1020 0 Vx1021 636.990790639369
Cx1020 x1020 xm1020 3.11541373257599e-14
Vx1020 xm1020 0 0
Gx1020_2 x1020 0 u2 0 -1.69697840920726e-07
Rx1021 x1021 0 1
Fxc1021_1020 x1021 0 Vx1020 -785.652076553797
Cx1021 x1021 xm1021 3.11541373257599e-14
Vx1021 xm1021 0 0
Gx1021_2 x1021 0 u2 0 0.000133323461106064
Rx1022 x1022 0 1
Fxc1022_1023 x1022 0 Vx1023 93.0625047322899
Cx1022 x1022 xm1022 1.22063164496342e-13
Vx1022 xm1022 0 0
Gx1022_2 x1022 0 u2 0 -5.03641784320086e-06
Rx1023 x1023 0 1
Fxc1023_1022 x1023 0 Vx1022 -359.175038648957
Cx1023 x1023 xm1023 1.22063164496342e-13
Vx1023 xm1023 0 0
Gx1023_2 x1023 0 u2 0 0.00180895557348396
Rx1024 x1024 0 1
Fxc1024_1025 x1024 0 Vx1025 224.107173585
Cx1024 x1024 xm1024 2.56056905033321e-14
Vx1024 xm1024 0 0
Gx1024_2 x1024 0 u2 0 -2.85141175082403e-08
Rx1025 x1025 0 1
Fxc1025_1024 x1025 0 Vx1024 -3342.58715214935
Cx1025 x1025 xm1025 2.56056905033321e-14
Vx1025 xm1025 0 0
Gx1025_2 x1025 0 u2 0 9.53109228379207e-05
Rx1026 x1026 0 1
Fxc1026_1027 x1026 0 Vx1027 2590.42388447807
Cx1026 x1026 xm1026 9.10350048138882e-15
Vx1026 xm1026 0 0
Gx1026_2 x1026 0 u2 0 -3.95670031491464e-09
Rx1027 x1027 0 1
Fxc1027_1026 x1027 0 Vx1026 -2400.8104179728
Cx1027 x1027 xm1027 9.10350048138882e-15
Vx1027 xm1027 0 0
Gx1027_2 x1027 0 u2 0 9.49928733684335e-06
Rx1028 x1028 0 1
Fxc1028_1029 x1028 0 Vx1029 1759.69003580951
Cx1028 x1028 xm1028 1.25795884003576e-14
Vx1028 xm1028 0 0
Gx1028_2 x1028 0 u2 0 -1.79311364661388e-08
Rx1029 x1029 0 1
Fxc1029_1028 x1029 0 Vx1028 -1774.47380035621
Cx1029 x1029 xm1029 1.25795884003576e-14
Vx1029 xm1029 0 0
Gx1029_2 x1029 0 u2 0 3.18183318697753e-05
Rx1030 x1030 0 1
Fxc1030_1031 x1030 0 Vx1031 8426.49482139967
Cx1030 x1030 xm1030 6.42832682389733e-15
Vx1030 xm1030 0 0
Gx1030_2 x1030 0 u2 0 -1.6810143794436e-09
Rx1031 x1031 0 1
Fxc1031_1030 x1031 0 Vx1030 -1457.02887146873
Cx1031 x1031 xm1031 6.42832682389733e-15
Vx1031 xm1031 0 0
Gx1031_2 x1031 0 u2 0 2.44928648420342e-06
Rx1032 x1032 0 1
Fxc1032_1033 x1032 0 Vx1033 178.427090061903
Cx1032 x1032 xm1032 3.78461462762688e-14
Vx1032 xm1032 0 0
Gx1032_2 x1032 0 u2 0 -5.01518715645875e-08
Rx1033 x1033 0 1
Fxc1033_1032 x1033 0 Vx1032 -2010.70047456672
Cx1033 x1033 xm1033 3.78461462762688e-14
Vx1033 xm1033 0 0
Gx1033_2 x1033 0 u2 0 0.000100840391955326
Rx1034 x1034 0 1
Fxc1034_1035 x1034 0 Vx1035 21256.1566440311
Cx1034 x1034 xm1034 7.47163154472276e-15
Vx1034 xm1034 0 0
Gx1034_2 x1034 0 u2 0 -1.35502392915902e-08
Rx1035 x1035 0 1
Fxc1035_1034 x1035 0 Vx1034 -422.660030061327
Cx1035 x1035 xm1035 7.47163154472277e-15
Vx1035 xm1035 0 0
Gx1035_2 x1035 0 u2 0 5.72714454632169e-06
Rx1036 x1036 0 1
Fxc1036_1037 x1036 0 Vx1037 2685.15989923165
Cx1036 x1036 xm1036 4.17550450563194e-14
Vx1036 xm1036 0 0
Gx1036_2 x1036 0 u2 0 -5.44628543455213e-07
Rx1037 x1037 0 1
Fxc1037_1036 x1037 0 Vx1036 -107.026435203432
Cx1037 x1037 xm1037 4.17550450563194e-14
Vx1037 xm1037 0 0
Gx1037_2 x1037 0 u2 0 5.82896515160487e-05
Rx1038 x1038 0 1
Fxc1038_1039 x1038 0 Vx1039 35759.404686904
Cx1038 x1038 xm1038 3.5696335326637e-13
Vx1038 xm1038 0 0
Gx1038_2 x1038 0 u2 0 -0.000195066100780617
Rx1039 x1039 0 1
Fxc1039_1038 x1039 0 Vx1038 -0.117841093405896
Cx1039 x1039 xm1039 3.5696335326637e-13
Vx1039 xm1039 0 0
Gx1039_2 x1039 0 u2 0 2.29868026024127e-05
Rx1040 x1040 0 1
Fxc1040_1041 x1040 0 Vx1041 782.940937910191
Cx1040 x1040 xm1040 1.92605907935797e-14
Vx1040 xm1040 0 0
Gx1040_2 x1040 0 u2 0 -1.90940090094287e-08
Rx1041 x1041 0 1
Fxc1041_1040 x1041 0 Vx1040 -1795.26563473352
Cx1041 x1041 xm1041 1.92605907935797e-14
Vx1041 xm1041 0 0
Gx1041_2 x1041 0 u2 0 3.42788182039197e-05
Rx1042 x1042 0 1
Fxc1042_1043 x1042 0 Vx1043 2083.12534858827
Cx1042 x1042 xm1042 4.96085474377487e-14
Vx1042 xm1042 0 0
Gx1042_2 x1042 0 u2 0 -4.09568525084372e-07
Rx1043 x1043 0 1
Fxc1043_1042 x1043 0 Vx1042 -102.151937604184
Cx1043 x1043 xm1043 4.96085474377487e-14
Vx1043 xm1043 0 0
Gx1043_2 x1043 0 u2 0 4.18382184190563e-05
Rx1044 x1044 0 1
Fxc1044_1045 x1044 0 Vx1045 4788.09370887249
Cx1044 x1044 xm1044 1.34382674878936e-14
Vx1044 xm1044 0 0
Gx1044_2 x1044 0 u2 0 -1.47424964305455e-08
Rx1045 x1045 0 1
Fxc1045_1044 x1045 0 Vx1044 -609.193085003472
Cx1045 x1045 xm1045 1.34382674878936e-14
Vx1045 xm1045 0 0
Gx1045_2 x1045 0 u2 0 8.98102688117667e-06
Rx1046 x1046 0 1
Fxc1046_1047 x1046 0 Vx1047 834.125771453118
Cx1046 x1046 xm1046 8.72908617003218e-15
Vx1046 xm1046 0 0
Gx1046_2 x1046 0 u2 0 -1.50517983676384e-09
Rx1047 x1047 0 1
Fxc1047_1046 x1047 0 Vx1046 -8404.38659087657
Cx1047 x1047 xm1047 8.72908617003218e-15
Vx1047 xm1047 0 0
Gx1047_2 x1047 0 u2 0 1.26501132369558e-05
Rx1048 x1048 0 1
Fxc1048_1049 x1048 0 Vx1049 774.542975989294
Cx1048 x1048 xm1048 1.41656257366965e-14
Vx1048 xm1048 0 0
Gx1048_2 x1048 0 u2 0 -4.74603290238197e-09
Rx1049 x1049 0 1
Fxc1049_1048 x1049 0 Vx1048 -3460.41173515052
Cx1049 x1049 xm1049 1.41656257366965e-14
Vx1049 xm1049 0 0
Gx1049_2 x1049 0 u2 0 1.64232279508131e-05
Rx1050 x1050 0 1
Fxc1050_1051 x1050 0 Vx1051 20.0706551775984
Cx1050 x1050 xm1050 6.46803689263805e-13
Vx1050 xm1050 0 0
Gx1050_2 x1050 0 u2 0 -0.000706517013427022
Rx1051 x1051 0 1
Fxc1051_1050 x1051 0 Vx1050 -69.0069944105614
Cx1051 x1051 xm1051 6.46803689263805e-13
Vx1051 xm1051 0 0
Gx1051_2 x1051 0 u2 0 0.048754615596525
Rx1052 x1052 0 1
Fxc1052_1053 x1052 0 Vx1053 98.4951815108806
Cx1052 x1052 xm1052 2.59067693849385e-14
Vx1052 xm1052 0 0
Gx1052_2 x1052 0 u2 0 -6.7061642317245e-09
Rx1053 x1053 0 1
Fxc1053_1052 x1053 0 Vx1052 -8204.09519742188
Cx1053 x1053 xm1053 2.59067693849385e-14
Vx1053 xm1053 0 0
Gx1053_2 x1053 0 u2 0 5.50180097666134e-05
Rx1054 x1054 0 1
Fxc1054_1055 x1054 0 Vx1055 16492.4068232391
Cx1054 x1054 xm1054 3.81925234457657e-15
Vx1054 xm1054 0 0
Gx1054_2 x1054 0 u2 0 -3.60216998452487e-09
Rx1055 x1055 0 1
Fxc1055_1054 x1055 0 Vx1054 -2277.16707417228
Cx1055 x1055 xm1055 3.81925234457657e-15
Vx1055 xm1055 0 0
Gx1055_2 x1055 0 u2 0 8.20274288433171e-06
Rx1056 x1056 0 1
Fxc1056_1057 x1056 0 Vx1057 140.156585829696
Cx1056 x1056 xm1056 5.61704850831073e-14
Vx1056 xm1056 0 0
Gx1056_2 x1056 0 u2 0 -2.50455204159313e-07
Rx1057 x1057 0 1
Fxc1057_1056 x1057 0 Vx1056 -1253.96234165531
Cx1057 x1057 xm1057 5.61704850831073e-14
Vx1057 xm1057 0 0
Gx1057_2 x1057 0 u2 0 0.000314061394287371
Rx1058 x1058 0 1
Fxc1058_1059 x1058 0 Vx1059 434.64479915759
Cx1058 x1058 xm1058 4.39028211648867e-14
Vx1058 xm1058 0 0
Gx1058_2 x1058 0 u2 0 -2.80851823913267e-07
Rx1059 x1059 0 1
Fxc1059_1058 x1059 0 Vx1058 -665.128856515029
Cx1059 x1059 xm1059 4.39028211648867e-14
Vx1059 xm1059 0 0
Gx1059_2 x1059 0 u2 0 0.000186802652489592
Rx1060 x1060 0 1
Fxc1060_1061 x1060 0 Vx1061 417.166158579639
Cx1060 x1060 xm1060 3.387890067806e-14
Vx1060 xm1060 0 0
Gx1060_2 x1060 0 u2 0 -9.06655850444836e-08
Rx1061 x1061 0 1
Fxc1061_1060 x1061 0 Vx1060 -1173.41145525554
Cx1061 x1061 xm1061 3.387890067806e-14
Vx1061 xm1061 0 0
Gx1061_2 x1061 0 u2 0 0.000106388036088642
Rx1062 x1062 0 1
Fxc1062_1063 x1062 0 Vx1063 12972.9182212671
Cx1062 x1062 xm1062 2.71987544670807e-14
Vx1062 xm1062 0 0
Gx1062_2 x1062 0 u2 0 -1.27674308226784e-07
Rx1063 x1063 0 1
Fxc1063_1062 x1063 0 Vx1062 -58.9467958658809
Cx1063 x1063 xm1063 2.71987544670807e-14
Vx1063 xm1063 0 0
Gx1063_2 x1063 0 u2 0 7.52599138436182e-06
Rx1064 x1064 0 1
Fxc1064_1065 x1064 0 Vx1065 93.1722462692019
Cx1064 x1064 xm1064 9.59156105724643e-14
Vx1064 xm1064 0 0
Gx1064_2 x1064 0 u2 0 -1.93796697261479e-06
Rx1065 x1065 0 1
Fxc1065_1064 x1065 0 Vx1064 -663.350902104362
Cx1065 x1065 xm1065 9.59156105724643e-14
Vx1065 xm1065 0 0
Gx1065_2 x1065 0 u2 0 0.00128555213953248
Rx1066 x1066 0 1
Fxc1066_1067 x1066 0 Vx1067 1556.15047288049
Cx1066 x1066 xm1066 2.29533381547327e-14
Vx1066 xm1066 0 0
Gx1066_2 x1066 0 u2 0 -1.50363920562097e-07
Rx1067 x1067 0 1
Fxc1067_1066 x1067 0 Vx1066 -697.148834537614
Cx1067 x1067 xm1067 2.29533381547327e-14
Vx1067 xm1067 0 0
Gx1067_2 x1067 0 u2 0 0.000104826031976372
Rx1068 x1068 0 1
Fxc1068_1069 x1068 0 Vx1069 5810.42639067816
Cx1068 x1068 xm1068 4.98360784941284e-15
Vx1068 xm1068 0 0
Gx1068_2 x1068 0 u2 0 -7.37758084731227e-09
Rx1069 x1069 0 1
Fxc1069_1068 x1069 0 Vx1068 -3967.37994612972
Cx1069 x1069 xm1069 4.98360784941284e-15
Vx1069 xm1069 0 0
Gx1069_2 x1069 0 u2 0 2.92696663045774e-05
Rx1070 x1070 0 1
Fxc1070_1071 x1070 0 Vx1071 3363.76840946582
Cx1070 x1070 xm1070 2.42570294480808e-15
Vx1070 xm1070 0 0
Gx1070_2 x1070 0 u2 0 -4.23437566670316e-10
Rx1071 x1071 0 1
Fxc1071_1070 x1071 0 Vx1070 -29365.5587054385
Cx1071 x1071 xm1071 2.42570294480808e-15
Vx1071 xm1071 0 0
Gx1071_2 x1071 0 u2 0 1.24344807221452e-05
Rx1072 x1072 0 1
Fxc1072_1073 x1072 0 Vx1073 15751.1714963422
Cx1072 x1072 xm1072 2.25473411609031e-15
Vx1072 xm1072 0 0
Gx1072_2 x1072 0 u2 0 -5.04902139546708e-10
Rx1073 x1073 0 1
Fxc1073_1072 x1073 0 Vx1072 -7308.923357827
Cx1073 x1073 xm1073 2.25473411609031e-15
Vx1073 xm1073 0 0
Gx1073_2 x1073 0 u2 0 3.69029104114976e-06
Rx1074 x1074 0 1
Fxc1074_1075 x1074 0 Vx1075 8.17108820913041
Cx1074 x1074 xm1074 1.48732812338964e-14
Vx1074 xm1074 0 0
Gx1074_2 x1074 0 u2 0 -8.33585658809323e-11
Rx1075 x1075 0 1
Fxc1075_1074 x1075 0 Vx1074 -326237.102318185
Cx1075 x1075 xm1075 1.48732812338964e-14
Vx1075 xm1075 0 0
Gx1075_2 x1075 0 u2 0 2.71946569863949e-05
Rx1076 x1076 0 1
Fxc1076_1077 x1076 0 Vx1077 21778.4890999364
Cx1076 x1076 xm1076 5.99616853581674e-15
Vx1076 xm1076 0 0
Gx1076_2 x1076 0 u2 0 -3.54677299850526e-09
Rx1077 x1077 0 1
Fxc1077_1076 x1077 0 Vx1076 -762.548916383372
Cx1077 x1077 xm1077 5.99616853581674e-15
Vx1077 xm1077 0 0
Gx1077_2 x1077 0 u2 0 2.70458790666799e-06
Rx1078 x1078 0 1
Fxc1078_1079 x1078 0 Vx1079 141.00851779169
Cx1078 x1078 xm1078 1.50857262477048e-14
Vx1078 xm1078 0 0
Gx1078_2 x1078 0 u2 0 -1.48609743012986e-09
Rx1079 x1079 0 1
Fxc1079_1078 x1079 0 Vx1078 -18781.9106907605
Cx1079 x1079 xm1079 1.50857262477048e-14
Vx1079 xm1079 0 0
Gx1079_2 x1079 0 u2 0 2.79117492104677e-05
Rx1080 x1080 0 1
Fxc1080_1081 x1080 0 Vx1081 1247.81479755534
Cx1080 x1080 xm1080 4.3895710802095e-15
Vx1080 xm1080 0 0
Gx1080_2 x1080 0 u2 0 -1.55258149106718e-10
Rx1081 x1081 0 1
Fxc1081_1080 x1081 0 Vx1080 -25216.8997130266
Cx1081 x1081 xm1081 4.3895710802095e-15
Vx1081 xm1081 0 0
Gx1081_2 x1081 0 u2 0 3.91512917565424e-06
Rx1082 x1082 0 1
Fxc1082_1083 x1082 0 Vx1083 510.542580925602
Cx1082 x1082 xm1082 1.55436740149653e-13
Vx1082 xm1082 0 0
Gx1082_2 x1082 0 u2 0 -7.20553871945691e-06
Rx1083 x1083 0 1
Fxc1083_1082 x1083 0 Vx1082 -49.9428567858924
Cx1083 x1083 xm1083 1.55436740149653e-13
Vx1083 xm1083 0 0
Gx1083_2 x1083 0 u2 0 0.000359865188331039
Rx1084 x1084 0 1
Fxc1084_1085 x1084 0 Vx1085 151024.665847056
Cx1084 x1084 xm1084 1.56758610576001e-15
Vx1084 xm1084 0 0
Gx1084_2 x1084 0 u2 0 -2.72472456814597e-10
Rx1085 x1085 0 1
Fxc1085_1084 x1085 0 Vx1084 -1651.23736791448
Cx1085 x1085 xm1085 1.56758610576001e-15
Vx1085 xm1085 0 0
Gx1085_2 x1085 0 u2 0 4.49916702419728e-07
Rx1086 x1086 0 1
Fxc1086_1087 x1086 0 Vx1087 163.02230726743
Cx1086 x1086 xm1086 3.97098834480777e-13
Vx1086 xm1086 0 0
Gx1086_2 x1086 0 u2 0 -0.000188366959888703
Rx1087 x1087 0 1
Fxc1087_1086 x1087 0 Vx1086 -24.9081790751194
Cx1087 x1087 xm1087 3.97098834480777e-13
Vx1087 xm1087 0 0
Gx1087_2 x1087 0 u2 0 0.00469187796874365
Rx1088 x1088 0 1
Fxc1088_1089 x1088 0 Vx1089 7274.04181818678
Cx1088 x1088 xm1088 1.20476536006176e-14
Vx1088 xm1088 0 0
Gx1088_2 x1088 0 u2 0 -1.41934430139079e-08
Rx1089 x1089 0 1
Fxc1089_1088 x1089 0 Vx1088 -583.950344752041
Cx1089 x1089 xm1089 1.20476536006176e-14
Vx1089 xm1089 0 0
Gx1089_2 x1089 0 u2 0 8.28826594118998e-06
Rx1090 x1090 0 1
Fxc1090_1091 x1090 0 Vx1091 1006621.6332794
Cx1090 x1090 xm1090 2.12416893515056e-16
Vx1090 xm1090 0 0
Gx1090_2 x1090 0 u2 0 -2.19899153692871e-10
Rx1091 x1091 0 1
Fxc1091_1090 x1091 0 Vx1090 -13829.8989283301
Cx1091 x1091 xm1091 2.12416893515056e-16
Vx1091 xm1091 0 0
Gx1091_2 x1091 0 u2 0 3.04118306999773e-06
Rx1092 x1092 0 1
Fxc1092_1093 x1092 0 Vx1093 330.013164620028
Cx1092 x1092 xm1092 9.7618575178155e-14
Vx1092 xm1092 0 0
Gx1092_2 x1092 0 u2 0 -1.62912393761235e-06
Rx1093 x1093 0 1
Fxc1093_1092 x1093 0 Vx1092 -200.350954663931
Cx1093 x1093 xm1093 9.7618575178155e-14
Vx1093 xm1093 0 0
Gx1093_2 x1093 0 u2 0 0.000326396536166495
Rx1094 x1094 0 1
Fxc1094_1095 x1094 0 Vx1095 133397.581862078
Cx1094 x1094 xm1094 1.87292384452854e-15
Vx1094 xm1094 0 0
Gx1094_2 x1094 0 u2 0 -1.07089827915982e-09
Rx1095 x1095 0 1
Fxc1095_1094 x1095 0 Vx1094 -1367.67399384489
Cx1095 x1095 xm1095 1.87292384452854e-15
Vx1095 xm1095 0 0
Gx1095_2 x1095 0 u2 0 1.46463972646013e-06
Rx1096 x1096 0 1
Fxc1096_1097 x1096 0 Vx1097 11718.6455399122
Cx1096 x1096 xm1096 1.43078355234661e-14
Vx1096 xm1096 0 0
Gx1096_2 x1096 0 u2 0 -6.4489324658816e-08
Rx1097 x1097 0 1
Fxc1097_1096 x1097 0 Vx1096 -266.753822570933
Cx1097 x1097 xm1097 1.43078355234661e-14
Vx1097 xm1097 0 0
Gx1097_2 x1097 0 u2 0 1.72027738677571e-05
Rx1098 x1098 0 1
Fxc1098_1099 x1098 0 Vx1099 123.206145027439
Cx1098 x1098 xm1098 1.25017605588615e-13
Vx1098 xm1098 0 0
Gx1098_2 x1098 0 u2 0 -3.89394270897075e-06
Rx1099 x1099 0 1
Fxc1099_1098 x1099 0 Vx1098 -375.436841285726
Cx1099 x1099 xm1099 1.25017605588615e-13
Vx1099 xm1099 0 0
Gx1099_2 x1099 0 u2 0 0.00146192955080356
Rx1100 x1100 0 1
Fxc1100_1101 x1100 0 Vx1101 604.016636842245
Cx1100 x1100 xm1100 2.53678675984263e-14
Vx1100 xm1100 0 0
Gx1100_2 x1100 0 u2 0 -3.40941350848639e-08
Rx1101 x1101 0 1
Fxc1101_1100 x1101 0 Vx1100 -1667.93702292329
Cx1101 x1101 xm1101 2.53678675984263e-14
Vx1101 xm1101 0 0
Gx1101_2 x1101 0 u2 0 5.68668701725924e-05
Rx1102 x1102 0 1
Fxc1102_1103 x1102 0 Vx1103 111170.077037626
Cx1102 x1102 xm1102 3.20804739778187e-16
Vx1102 xm1102 0 0
Gx1102_2 x1102 0 u2 0 -2.8598027721088e-10
Rx1103 x1103 0 1
Fxc1103_1102 x1103 0 Vx1102 -56926.011169663
Cx1103 x1103 xm1103 3.20804739778187e-16
Vx1103 xm1103 0 0
Gx1103_2 x1103 0 u2 0 1.62797164548099e-05
Rx1104 x1104 0 1
Fxc1104_1105 x1104 0 Vx1105 4859.24738828328
Cx1104 x1104 xm1104 2.27190048287476e-14
Vx1104 xm1104 0 0
Gx1104_2 x1104 0 u2 0 -3.55382368479671e-08
Rx1105 x1105 0 1
Fxc1105_1104 x1105 0 Vx1104 -262.368118108764
Cx1105 x1105 xm1105 2.27190048287476e-14
Vx1105 xm1105 0 0
Gx1105_2 x1105 0 u2 0 9.32410032270466e-06
Rx1106 x1106 0 1
Fxc1106_1107 x1106 0 Vx1107 104.508606374775
Cx1106 x1106 xm1106 2.2084230164543e-13
Vx1106 xm1106 0 0
Gx1106_2 x1106 0 u2 0 -2.57365176405953e-05
Rx1107 x1107 0 1
Fxc1107_1106 x1107 0 Vx1106 -132.849612747434
Cx1107 x1107 xm1107 2.2084230164543e-13
Vx1107 xm1107 0 0
Gx1107_2 x1107 0 u2 0 0.00341908640202058
Rx1108 x1108 0 1
Fxc1108_1109 x1108 0 Vx1109 2371.90945245139
Cx1108 x1108 xm1108 2.43012562210102e-13
Vx1108 xm1108 0 0
Gx1108_2 x1108 0 u2 0 -4.48179009037208e-05
Rx1109 x1109 0 1
Fxc1109_1108 x1109 0 Vx1108 -4.94009074476777
Cx1109 x1109 xm1109 2.43012562210102e-13
Vx1109 xm1109 0 0
Gx1109_2 x1109 0 u2 0 0.00022140449745439
Rx1110 x1110 0 1
Fxc1110_1111 x1110 0 Vx1111 691.601335650312
Cx1110 x1110 xm1110 3.92393390132605e-14
Vx1110 xm1110 0 0
Gx1110_2 x1110 0 u2 0 -1.16654081192051e-07
Rx1111 x1111 0 1
Fxc1111_1110 x1111 0 Vx1110 -635.538481425168
Cx1111 x1111 xm1111 3.92393390132605e-14
Vx1111 xm1111 0 0
Gx1111_2 x1111 0 u2 0 7.41381576128444e-05
Rx1112 x1112 0 1
Fxc1112_1113 x1112 0 Vx1113 159.360437536608
Cx1112 x1112 xm1112 2.14454644620413e-14
Vx1112 xm1112 0 0
Gx1112_2 x1112 0 u2 0 -5.45709752429576e-09
Rx1113 x1113 0 1
Fxc1113_1112 x1113 0 Vx1112 -9133.48198095708
Cx1113 x1113 xm1113 2.14454644620413e-14
Vx1113 xm1113 0 0
Gx1113_2 x1113 0 u2 0 4.98423019064809e-05
Rx1114 x1114 0 1
Fxc1114_1115 x1114 0 Vx1115 199.640214060821
Cx1114 x1114 xm1114 3.69189637458766e-14
Vx1114 xm1114 0 0
Gx1114_2 x1114 0 u2 0 -3.77140196638512e-08
Rx1115 x1115 0 1
Fxc1115_1114 x1115 0 Vx1114 -2530.17947034386
Cx1115 x1115 xm1115 3.69189637458766e-14
Vx1115 xm1115 0 0
Gx1115_2 x1115 0 u2 0 9.54232382976209e-05
Rx1116 x1116 0 1
Fxc1116_1117 x1116 0 Vx1117 491.300797636117
Cx1116 x1116 xm1116 1.78601578922452e-14
Vx1116 xm1116 0 0
Gx1116_2 x1116 0 u2 0 -7.52067955417449e-09
Rx1117 x1117 0 1
Fxc1117_1116 x1117 0 Vx1116 -4524.82741365591
Cx1117 x1117 xm1117 1.78601578922452e-14
Vx1117 xm1117 0 0
Gx1117_2 x1117 0 u2 0 3.40297770160503e-05
Rx1118 x1118 0 1
Fxc1118_1119 x1118 0 Vx1119 26713.3341699692
Cx1118 x1118 xm1118 3.02453155184689e-14
Vx1118 xm1118 0 0
Gx1118_2 x1118 0 u2 0 -6.81879850847876e-08
Rx1119 x1119 0 1
Fxc1119_1118 x1119 0 Vx1118 -28.4189281794892
Cx1119 x1119 xm1119 3.02453155184689e-14
Vx1119 xm1119 0 0
Gx1119_2 x1119 0 u2 0 1.93782945082866e-06
Rx1120 x1120 0 1
Fxc1120_1121 x1120 0 Vx1121 493.560269581913
Cx1120 x1120 xm1120 3.68500092864944e-14
Vx1120 xm1120 0 0
Gx1120_2 x1120 0 u2 0 -7.43673004312087e-08
Rx1121 x1121 0 1
Fxc1121_1120 x1121 0 Vx1120 -1067.61389635874
Cx1121 x1121 xm1121 3.68500092864944e-14
Vx1121 xm1121 0 0
Gx1121_2 x1121 0 u2 0 7.93955633750437e-05
Rx1122 x1122 0 1
Fxc1122_1123 x1122 0 Vx1123 393.045587075839
Cx1122 x1122 xm1122 4.62675941996372e-14
Vx1122 xm1122 0 0
Gx1122_2 x1122 0 u2 0 -1.39998439399693e-07
Rx1123 x1123 0 1
Fxc1123_1122 x1123 0 Vx1122 -789.161372956843
Cx1123 x1123 xm1123 4.62675941996372e-14
Vx1123 xm1123 0 0
Gx1123_2 x1123 0 u2 0 0.000110481360648477
Rx1124 x1124 0 1
Fxc1124_1125 x1124 0 Vx1125 1045.5285113103
Cx1124 x1124 xm1124 2.94176684113735e-15
Vx1124 xm1124 0 0
Gx1124_2 x1124 0 u2 0 -1.62887517186097e-10
Rx1125 x1125 0 1
Fxc1125_1124 x1125 0 Vx1124 -77621.6648129607
Cx1125 x1125 xm1125 2.94176684113735e-15
Vx1125 xm1125 0 0
Gx1125_2 x1125 0 u2 0 1.26436002612346e-05
Rx1126 x1126 0 1
Fxc1126_1127 x1126 0 Vx1127 5658.19332327565
Cx1126 x1126 xm1126 9.26868572070505e-15
Vx1126 xm1126 0 0
Gx1126_2 x1126 0 u2 0 -6.96188178670615e-09
Rx1127 x1127 0 1
Fxc1127_1126 x1127 0 Vx1126 -1544.38197378395
Cx1127 x1127 xm1127 9.26868572070505e-15
Vx1127 xm1127 0 0
Gx1127_2 x1127 0 u2 0 1.07518047350038e-05
Rx1128 x1128 0 1
Fxc1128_1129 x1128 0 Vx1129 366.451608395772
Cx1128 x1128 xm1128 4.05009397042418e-14
Vx1128 xm1128 0 0
Gx1128_2 x1128 0 u2 0 -5.38528331460671e-08
Rx1129 x1129 0 1
Fxc1129_1128 x1129 0 Vx1128 -1236.43706462843
Cx1129 x1129 xm1129 4.05009397042418e-14
Vx1129 xm1129 0 0
Gx1129_2 x1129 0 u2 0 6.65856389370479e-05
Rx1130 x1130 0 1
Fxc1130_1131 x1130 0 Vx1131 1427.82729202391
Cx1130 x1130 xm1130 4.03994326186591e-15
Vx1130 xm1130 0 0
Gx1130_2 x1130 0 u2 0 -4.45138029836028e-10
Rx1131 x1131 0 1
Fxc1131_1130 x1131 0 Vx1130 -31602.700632607
Cx1131 x1131 xm1131 4.03994326186591e-15
Vx1131 xm1131 0 0
Gx1131_2 x1131 0 u2 0 1.40675638970965e-05
Rx1132 x1132 0 1
Fxc1132_1133 x1132 0 Vx1133 8319.79745095293
Cx1132 x1132 xm1132 1.4939511468885e-13
Vx1132 xm1132 0 0
Gx1132_2 x1132 0 u2 0 -1.13039380404279e-05
Rx1133 x1133 0 1
Fxc1133_1132 x1133 0 Vx1132 -3.91423466532942
Cx1133 x1133 xm1133 1.4939511468885e-13
Vx1133 xm1133 0 0
Gx1133_2 x1133 0 u2 0 4.42462661325786e-05
Rx1134 x1134 0 1
Fxc1134_1135 x1134 0 Vx1135 11538.8025427113
Cx1134 x1134 xm1134 1.24148427126151e-14
Vx1134 xm1134 0 0
Gx1134_2 x1134 0 u2 0 -3.61437428492281e-09
Rx1135 x1135 0 1
Fxc1135_1134 x1135 0 Vx1134 -408.202926156697
Cx1135 x1135 xm1135 1.24148427126152e-14
Vx1135 xm1135 0 0
Gx1135_2 x1135 0 u2 0 1.47539815933101e-06
Rx1136 x1136 0 1
Fxc1136_1137 x1136 0 Vx1137 356.545057646723
Cx1136 x1136 xm1136 3.04285853351407e-14
Vx1136 xm1136 0 0
Gx1136_2 x1136 0 u2 0 -2.76830164562241e-08
Rx1137 x1137 0 1
Fxc1137_1136 x1137 0 Vx1136 -2297.66108339779
Cx1137 x1137 xm1137 3.04285853351407e-14
Vx1137 xm1137 0 0
Gx1137_2 x1137 0 u2 0 6.36061895825267e-05
Rx1138 x1138 0 1
Fxc1138_1139 x1138 0 Vx1139 149564.131055872
Cx1138 x1138 xm1138 2.80028892882111e-16
Vx1138 xm1138 0 0
Gx1138_2 x1138 0 u2 0 -7.65769422751694e-11
Rx1139 x1139 0 1
Fxc1139_1138 x1139 0 Vx1138 -65558.8490641051
Cx1139 x1139 xm1139 2.80028892882111e-16
Vx1139 xm1139 0 0
Gx1139_2 x1139 0 u2 0 5.02029620040852e-06
Rx1140 x1140 0 1
Fxc1140_1141 x1140 0 Vx1141 893.590212536684
Cx1140 x1140 xm1140 5.53119643557016e-15
Vx1140 xm1140 0 0
Gx1140_2 x1140 0 u2 0 -5.94999100285696e-10
Rx1141 x1141 0 1
Fxc1141_1140 x1141 0 Vx1140 -28697.3977506826
Cx1141 x1141 xm1141 5.53119643557016e-15
Vx1141 xm1141 0 0
Gx1141_2 x1141 0 u2 0 1.70749258421969e-05
Rx1142 x1142 0 1
Fxc1142_1143 x1142 0 Vx1143 18179.6527795021
Cx1142 x1142 xm1142 3.62906157244733e-15
Vx1142 xm1142 0 0
Gx1142_2 x1142 0 u2 0 -7.25901929981006e-10
Rx1143 x1143 0 1
Fxc1143_1142 x1143 0 Vx1142 -3240.85099700554
Cx1143 x1143 xm1143 3.62906157244733e-15
Vx1143 xm1143 0 0
Gx1143_2 x1143 0 u2 0 2.35253999350719e-06
Rx1144 x1144 0 1
Fxc1144_1145 x1144 0 Vx1145 958.269077504141
Cx1144 x1144 xm1144 2.43563137386751e-14
Vx1144 xm1144 0 0
Gx1144_2 x1144 0 u2 0 -1.8878445149944e-08
Rx1145 x1145 0 1
Fxc1145_1144 x1145 0 Vx1144 -1402.31900722099
Cx1145 x1145 xm1145 2.43563137386751e-14
Vx1145 xm1145 0 0
Gx1145_2 x1145 0 u2 0 2.64736024605454e-05
Rx1146 x1146 0 1
Fxc1146_1147 x1146 0 Vx1147 8041.95900577969
Cx1146 x1146 xm1146 7.64511008833615e-15
Vx1146 xm1146 0 0
Gx1146_2 x1146 0 u2 0 -2.63290758008851e-09
Rx1147 x1147 0 1
Fxc1147_1146 x1147 0 Vx1146 -1685.81863067129
Cx1147 x1147 xm1147 7.64511008833615e-15
Vx1147 xm1147 0 0
Gx1147_2 x1147 0 u2 0 4.43860465134888e-06
Rx1148 x1148 0 1
Fxc1148_1149 x1148 0 Vx1149 824.974373147359
Cx1148 x1148 xm1148 3.31932360252982e-14
Vx1148 xm1148 0 0
Gx1148_2 x1148 0 u2 0 -7.64638362102977e-08
Rx1149 x1149 0 1
Fxc1149_1148 x1149 0 Vx1148 -830.8972290859
Cx1149 x1149 xm1149 3.31932360252982e-14
Vx1149 xm1149 0 0
Gx1149_2 x1149 0 u2 0 6.35335896324145e-05
Rx1150 x1150 0 1
Fxc1150_1151 x1150 0 Vx1151 39.8478517389542
Cx1150 x1150 xm1150 3.91990471759038e-13
Vx1150 xm1150 0 0
Gx1150_2 x1150 0 u2 0 -0.000176163857726359
Rx1151 x1151 0 1
Fxc1151_1150 x1151 0 Vx1150 -135.643395145431
Cx1151 x1151 xm1151 3.91990471759038e-13
Vx1151 xm1151 0 0
Gx1151_2 x1151 0 u2 0 0.02389546376392
Rx1152 x1152 0 1
Fxc1152_1153 x1152 0 Vx1153 7415.8466967697
Cx1152 x1152 xm1152 1.62720964829041e-14
Vx1152 xm1152 0 0
Gx1152_2 x1152 0 u2 0 -3.24848887586088e-08
Rx1153 x1153 0 1
Fxc1153_1152 x1153 0 Vx1152 -410.061245643613
Cx1153 x1153 xm1153 1.62720964829041e-14
Vx1153 xm1153 0 0
Gx1153_2 x1153 0 u2 0 1.33207939489493e-05
Rx1154 x1154 0 1
Fxc1154_1155 x1154 0 Vx1155 550.54521148892
Cx1154 x1154 xm1154 8.80522494224567e-14
Vx1154 xm1154 0 0
Gx1154_2 x1154 0 u2 0 -1.16597747495329e-06
Rx1155 x1155 0 1
Fxc1155_1154 x1155 0 Vx1154 -188.777966798872
Cx1155 x1155 xm1155 8.80522494224567e-14
Vx1155 xm1155 0 0
Gx1155_2 x1155 0 u2 0 0.000220110857054964
Rx1156 x1156 0 1
Fxc1156_1157 x1156 0 Vx1157 4.18409898701301
Cx1156 x1156 xm1156 7.67229662280685e-13
Vx1156 xm1156 0 0
Gx1156_2 x1156 0 u2 0 -0.000233899439118769
Rx1157 x1157 0 1
Fxc1157_1156 x1157 0 Vx1156 -365.781574536642
Cx1157 x1157 xm1157 7.67229662280685e-13
Vx1157 xm1157 0 0
Gx1157_2 x1157 0 u2 0 0.0855561051241005
Rx1158 x1158 0 1
Fxc1158_1159 x1158 0 Vx1159 1.53910429470818
Cx1158 x1158 xm1158 4.92776735733474e-13
Vx1158 xm1158 0 0
Gx1158_2 x1158 0 u2 0 -2.31139972137463e-05
Rx1159 x1159 0 1
Fxc1159_1158 x1159 0 Vx1158 -2236.91020350738
Cx1159 x1159 xm1159 4.92776735733474e-13
Vx1159 xm1159 0 0
Gx1159_2 x1159 0 u2 0 0.0517039362112704
Rx1160 x1160 0 1
Fxc1160_1161 x1160 0 Vx1161 150.854880601286
Cx1160 x1160 xm1160 1.65994637491899e-14
Vx1160 xm1160 0 0
Gx1160_2 x1160 0 u2 0 -1.63907804610197e-09
Rx1161 x1161 0 1
Fxc1161_1160 x1161 0 Vx1160 -19677.8823066489
Cx1161 x1161 xm1161 1.65994637491899e-14
Vx1161 xm1161 0 0
Gx1161_2 x1161 0 u2 0 3.22535848826065e-05
Rx1162 x1162 0 1
Fxc1162_1163 x1162 0 Vx1163 5973.69894274732
Cx1162 x1162 xm1162 1.52443737477815e-14
Vx1162 xm1162 0 0
Gx1162_2 x1162 0 u2 0 -7.16640749180273e-09
Rx1163 x1163 0 1
Fxc1163_1162 x1163 0 Vx1162 -594.589237404974
Cx1163 x1163 xm1163 1.52443737477815e-14
Vx1163 xm1163 0 0
Gx1163_2 x1163 0 u2 0 4.26106876548428e-06
Rx1164 x1164 0 1
Fxc1164_1165 x1164 0 Vx1165 111.683148228054
Cx1164 x1164 xm1164 2.73296090832205e-13
Vx1164 xm1164 0 0
Gx1164_2 x1164 0 u2 0 -3.88020230081831e-05
Rx1165 x1165 0 1
Fxc1165_1164 x1165 0 Vx1164 -109.883108235608
Cx1165 x1165 xm1165 2.73296090832205e-13
Vx1165 xm1165 0 0
Gx1165_2 x1165 0 u2 0 0.00426368689396875
Rx1166 x1166 0 1
Fxc1166_1167 x1166 0 Vx1167 529.191521623437
Cx1166 x1166 xm1166 2.87228473774017e-14
Vx1166 xm1166 0 0
Gx1166_2 x1166 0 u2 0 -2.05656287133461e-08
Rx1167 x1167 0 1
Fxc1167_1166 x1167 0 Vx1166 -1924.67650373784
Cx1167 x1167 xm1167 2.87228473774017e-14
Vx1167 xm1167 0 0
Gx1167_2 x1167 0 u2 0 3.95821823691733e-05
Rx1168 x1168 0 1
Fxc1168_1169 x1168 0 Vx1169 1163.47534613422
Cx1168 x1168 xm1168 4.66685567425351e-14
Vx1168 xm1168 0 0
Gx1168_2 x1168 0 u2 0 -1.28378315978994e-07
Rx1169 x1169 0 1
Fxc1169_1168 x1169 0 Vx1168 -336.17165522018
Cx1169 x1169 xm1169 4.66685567425351e-14
Vx1169 xm1169 0 0
Gx1169_2 x1169 0 u2 0 4.31571509770376e-05
Rx1170 x1170 0 1
Fxc1170_1171 x1170 0 Vx1171 710.163903512532
Cx1170 x1170 xm1170 5.7196013910315e-14
Vx1170 xm1170 0 0
Gx1170_2 x1170 0 u2 0 -2.22014488780856e-07
Rx1171 x1171 0 1
Fxc1171_1170 x1171 0 Vx1170 -369.536285734102
Cx1171 x1171 xm1171 5.7196013910315e-14
Vx1171 xm1171 0 0
Gx1171_2 x1171 0 u2 0 8.20424095632329e-05
Rx1172 x1172 0 1
Fxc1172_1173 x1172 0 Vx1173 193.630058649167
Cx1172 x1172 xm1172 1.75688323351063e-13
Vx1172 xm1172 0 0
Gx1172_2 x1172 0 u2 0 -1.12709789894303e-05
Rx1173 x1173 0 1
Fxc1173_1172 x1173 0 Vx1172 -148.408819666664
Cx1173 x1173 xm1173 1.75688323351063e-13
Vx1173 xm1173 0 0
Gx1173_2 x1173 0 u2 0 0.00167271268830912
Rx1174 x1174 0 1
Fxc1174_1175 x1174 0 Vx1175 12954.0722479593
Cx1174 x1174 xm1174 6.22004467114814e-14
Vx1174 xm1174 0 0
Gx1174_2 x1174 0 u2 0 -4.10682077129726e-07
Rx1175 x1175 0 1
Fxc1175_1174 x1175 0 Vx1174 -17.857611576843
Cx1175 x1175 xm1175 6.22004467114814e-14
Vx1175 xm1175 0 0
Gx1175_2 x1175 0 u2 0 7.33380101495373e-06
Rx1176 x1176 0 1
Fxc1176_1177 x1176 0 Vx1177 14271.5171680843
Cx1176 x1176 xm1176 1.41434995567386e-14
Vx1176 xm1176 0 0
Gx1176_2 x1176 0 u2 0 -1.14932194987322e-08
Rx1177 x1177 0 1
Fxc1177_1176 x1177 0 Vx1176 -305.233090503257
Cx1177 x1177 xm1177 1.41434995567386e-14
Vx1177 xm1177 0 0
Gx1177_2 x1177 0 u2 0 3.50811090743032e-06
Rx1178 x1178 0 1
Fxc1178_1179 x1178 0 Vx1179 323.712329039208
Cx1178 x1178 xm1178 5.26768043602151e-14
Vx1178 xm1178 0 0
Gx1178_2 x1178 0 u2 0 -1.38786097811487e-07
Rx1179 x1179 0 1
Fxc1179_1178 x1179 0 Vx1178 -980.937248756173
Cx1179 x1179 xm1179 5.26768043602151e-14
Vx1179 xm1179 0 0
Gx1179_2 x1179 0 u2 0 0.000136140452952805
Rx1180 x1180 0 1
Fxc1180_1181 x1180 0 Vx1181 1343.6184633664
Cx1180 x1180 xm1180 5.31047753536345e-14
Vx1180 xm1180 0 0
Gx1180_2 x1180 0 u2 0 -2.02023760407565e-07
Rx1181 x1181 0 1
Fxc1181_1180 x1181 0 Vx1180 -240.120308883562
Cx1181 x1181 xm1181 5.31047753536345e-14
Vx1181 xm1181 0 0
Gx1181_2 x1181 0 u2 0 4.85100077508831e-05
Rx1182 x1182 0 1
Fxc1182_1183 x1182 0 Vx1183 761.782081126751
Cx1182 x1182 xm1182 1.32036835764334e-14
Vx1182 xm1182 0 0
Gx1182_2 x1182 0 u2 0 -1.70657221221085e-09
Rx1183 x1183 0 1
Fxc1183_1182 x1183 0 Vx1182 -6932.28810890847
Cx1183 x1183 xm1183 1.32036835764334e-14
Vx1183 xm1183 0 0
Gx1183_2 x1183 0 u2 0 1.18304502537029e-05
Rx1184 x1184 0 1
Fxc1184_1185 x1184 0 Vx1185 40.0238746952908
Cx1184 x1184 xm1184 5.7822019650203e-13
Vx1184 xm1184 0 0
Gx1184_2 x1184 0 u2 0 -0.00047278801294426
Rx1185 x1185 0 1
Fxc1185_1184 x1185 0 Vx1184 -73.29653304629
Cx1185 x1185 xm1185 5.7822019650203e-13
Vx1185 xm1185 0 0
Gx1185_2 x1185 0 u2 0 0.0346537222146587
Rx1186 x1186 0 1
Fxc1186_1187 x1186 0 Vx1187 674.777596183298
Cx1186 x1186 xm1186 1.02035760349352e-13
Vx1186 xm1186 0 0
Gx1186_2 x1186 0 u2 0 -1.09109373300298e-06
Rx1187 x1187 0 1
Fxc1187_1186 x1187 0 Vx1186 -132.796787785316
Cx1187 x1187 xm1187 1.02035760349352e-13
Vx1187 xm1187 0 0
Gx1187_2 x1187 0 u2 0 0.000144893742915486
Rx1188 x1188 0 1
Fxc1188_1189 x1188 0 Vx1189 18108.0876442907
Cx1188 x1188 xm1188 2.40247346728811e-14
Vx1188 xm1188 0 0
Gx1188_2 x1188 0 u2 0 -3.98238152048716e-08
Rx1189 x1189 0 1
Fxc1189_1188 x1189 0 Vx1188 -90.1600647626225
Cx1189 x1189 xm1189 2.40247346728811e-14
Vx1189 xm1189 0 0
Gx1189_2 x1189 0 u2 0 3.59051775796594e-06
Rx1190 x1190 0 1
Fxc1190_1191 x1190 0 Vx1191 154.955738781269
Cx1190 x1190 xm1190 3.08852421707331e-14
Vx1190 xm1190 0 0
Gx1190_2 x1190 0 u2 0 -6.80692513851505e-09
Rx1191 x1191 0 1
Fxc1191_1190 x1191 0 Vx1190 -6436.53634941262
Cx1191 x1191 xm1191 3.08852421707331e-14
Vx1191 xm1191 0 0
Gx1191_2 x1191 0 u2 0 4.38130210817826e-05
Rx1192 x1192 0 1
Fxc1192_1193 x1192 0 Vx1193 1522.74713931895
Cx1192 x1192 xm1192 1.63019845419542e-14
Vx1192 xm1192 0 0
Gx1192_2 x1192 0 u2 0 -7.26392412791558e-09
Rx1193 x1193 0 1
Fxc1193_1192 x1193 0 Vx1192 -2366.83097721828
Cx1193 x1193 xm1193 1.63019845419542e-14
Vx1193 xm1193 0 0
Gx1193_2 x1193 0 u2 0 1.71924806421139e-05
Rx1194 x1194 0 1
Fxc1194_1195 x1194 0 Vx1195 110.537515069427
Cx1194 x1194 xm1194 6.41736383827721e-13
Vx1194 xm1194 0 0
Gx1194_2 x1194 0 u2 0 -0.00061333543240601
Rx1195 x1195 0 1
Fxc1195_1194 x1195 0 Vx1194 -23.0420317221486
Cx1195 x1195 xm1195 6.41736383827721e-13
Vx1195 xm1195 0 0
Gx1195_2 x1195 0 u2 0 0.014132494489817
Rx1196 x1196 0 1
Fxc1196_1197 x1196 0 Vx1197 24.960665570798
Cx1196 x1196 xm1196 2.85479875469681e-14
Vx1196 xm1196 0 0
Gx1196_2 x1196 0 u2 0 -9.70040035585148e-10
Rx1197 x1197 0 1
Fxc1197_1196 x1197 0 Vx1196 -47648.3923878378
Cx1197 x1197 xm1197 2.85479875469681e-14
Vx1197 xm1197 0 0
Gx1197_2 x1197 0 u2 0 4.62208482474732e-05
Rx1198 x1198 0 1
Fxc1198_1199 x1198 0 Vx1199 29.6943581226018
Cx1198 x1198 xm1198 5.3285703820123e-13
Vx1198 xm1198 0 0
Gx1198_2 x1198 0 u2 0 -0.000368693356736194
Rx1199 x1199 0 1
Fxc1199_1198 x1199 0 Vx1198 -120.002011248125
Cx1199 x1199 xm1199 5.3285703820123e-13
Vx1199 xm1199 0 0
Gx1199_2 x1199 0 u2 0 0.0442439443421656
Rx1200 x1200 0 1
Fxc1200_1201 x1200 0 Vx1201 245.108620915453
Cx1200 x1200 xm1200 3.03498701128083e-14
Vx1200 xm1200 0 0
Gx1200_2 x1200 0 u2 0 -9.02545440456516e-09
Rx1201 x1201 0 1
Fxc1201_1200 x1201 0 Vx1200 -4320.47233343833
Cx1201 x1201 xm1201 3.03498701128083e-14
Vx1201 xm1201 0 0
Gx1201_2 x1201 0 u2 0 3.89942260516329e-05
Rx1202 x1202 0 1
Fxc1202_1203 x1202 0 Vx1203 537.250528482313
Cx1202 x1202 xm1202 1.01462685758652e-13
Vx1202 xm1202 0 0
Gx1202_2 x1202 0 u2 0 -1.3768609761927e-06
Rx1203 x1203 0 1
Fxc1203_1202 x1203 0 Vx1202 -180.100871356267
Cx1203 x1203 xm1203 1.01462685758652e-13
Vx1203 xm1203 0 0
Gx1203_2 x1203 0 u2 0 0.000247973861548745
Rx1204 x1204 0 1
Fxc1204_1205 x1204 0 Vx1205 1176.72327136142
Cx1204 x1204 xm1204 1.02325988713972e-13
Vx1204 xm1204 0 0
Gx1204_2 x1204 0 u2 0 -1.68807511588321e-06
Rx1205 x1205 0 1
Fxc1205_1204 x1205 0 Vx1204 -81.6533117941909
Cx1205 x1205 xm1205 1.02325988713972e-13
Vx1205 xm1205 0 0
Gx1205_2 x1205 0 u2 0 0.000137836923769227
Rx1206 x1206 0 1
Fxc1206_1207 x1206 0 Vx1207 77.7622993065366
Cx1206 x1206 xm1206 1.41000112840634e-13
Vx1206 xm1206 0 0
Gx1206_2 x1206 0 u2 0 -2.63169478471067e-06
Rx1207 x1207 0 1
Fxc1207_1206 x1207 0 Vx1206 -736.709104997434
Cx1207 x1207 xm1207 1.41000112840634e-13
Vx1207 xm1207 0 0
Gx1207_2 x1207 0 u2 0 0.00193879350947061
Rx1208 x1208 0 1
Fxc1208_1209 x1208 0 Vx1209 199.532511128906
Cx1208 x1208 xm1208 1.32754836741219e-13
Vx1208 xm1208 0 0
Gx1208_2 x1208 0 u2 0 -1.70470170027686e-06
Rx1209 x1209 0 1
Fxc1209_1208 x1209 0 Vx1208 -291.326969437204
Cx1209 x1209 xm1209 1.32754836741219e-13
Vx1209 xm1209 0 0
Gx1209_2 x1209 0 u2 0 0.000496625580136107
Rx1210 x1210 0 1
Fxc1210_1211 x1210 0 Vx1211 516.246460573248
Cx1210 x1210 xm1210 1.26702180135926e-14
Vx1210 xm1210 0 0
Gx1210_2 x1210 0 u2 0 -9.31662898765873e-10
Rx1211 x1211 0 1
Fxc1211_1210 x1211 0 Vx1210 -13559.6066155356
Cx1211 x1211 xm1211 1.26702180135926e-14
Vx1211 xm1211 0 0
Gx1211_2 x1211 0 u2 0 1.26329824055548e-05
Rx1212 x1212 0 1
Fxc1212_1213 x1212 0 Vx1213 469.841654279092
Cx1212 x1212 xm1212 3.01789464736231e-14
Vx1212 xm1212 0 0
Gx1212_2 x1212 0 u2 0 -9.49112064934095e-09
Rx1213 x1213 0 1
Fxc1213_1212 x1213 0 Vx1212 -2482.57470102622
Cx1213 x1213 xm1213 3.01789464736231e-14
Vx1213 xm1213 0 0
Gx1213_2 x1213 0 u2 0 2.35624160084414e-05
Rx1214 x1214 0 1
Fxc1214_1215 x1214 0 Vx1215 487.563238195966
Cx1214 x1214 xm1214 9.70484385291882e-14
Vx1214 xm1214 0 0
Gx1214_2 x1214 0 u2 0 -9.97124057591693e-07
Rx1215 x1215 0 1
Fxc1215_1214 x1215 0 Vx1214 -238.362281502606
Cx1215 x1215 xm1215 9.70484385291883e-14
Vx1215 xm1215 0 0
Gx1215_2 x1215 0 u2 0 0.000237676765308691
Rx1216 x1216 0 1
Fxc1216_1217 x1216 0 Vx1217 788.132449380105
Cx1216 x1216 xm1216 3.43607207471199e-14
Vx1216 xm1216 0 0
Gx1216_2 x1216 0 u2 0 -3.19335635523789e-08
Rx1217 x1217 0 1
Fxc1217_1216 x1217 0 Vx1216 -1133.69551966872
Cx1217 x1217 xm1217 3.43607207471199e-14
Vx1217 xm1217 0 0
Gx1217_2 x1217 0 u2 0 3.62029379263883e-05
Rx1218 x1218 0 1
Fxc1218_1219 x1218 0 Vx1219 276.431040299342
Cx1218 x1218 xm1218 1.54871227469822e-13
Vx1218 xm1218 0 0
Gx1218_2 x1218 0 u2 0 -4.55953889285e-06
Rx1219 x1219 0 1
Fxc1219_1218 x1219 0 Vx1218 -165.930800413054
Cx1219 x1219 xm1219 1.54871227469822e-13
Vx1219 xm1219 0 0
Gx1219_2 x1219 0 u2 0 0.000756567938005048
Rx1220 x1220 0 1
Fxc1220_1221 x1220 0 Vx1221 170.452686566085
Cx1220 x1220 xm1220 6.44307967443506e-14
Vx1220 xm1220 0 0
Gx1220_2 x1220 0 u2 0 -6.48430654140735e-08
Rx1221 x1221 0 1
Fxc1221_1220 x1221 0 Vx1220 -1529.13848831447
Cx1221 x1221 xm1221 6.44307967443506e-14
Vx1221 xm1221 0 0
Gx1221_2 x1221 0 u2 0 9.91540270249528e-05
Rx1222 x1222 0 1
Fxc1222_1223 x1222 0 Vx1223 9145.70669848558
Cx1222 x1222 xm1222 2.24357038343354e-14
Vx1222 xm1222 0 0
Gx1222_2 x1222 0 u2 0 -2.48068321412333e-08
Rx1223 x1223 0 1
Fxc1223_1222 x1223 0 Vx1222 -238.737602518704
Cx1223 x1223 xm1223 2.24357038343354e-14
Vx1223 xm1223 0 0
Gx1223_2 x1223 0 u2 0 5.92232363148196e-06
Rx1224 x1224 0 1
Fxc1224_1225 x1224 0 Vx1225 1687.70634504343
Cx1224 x1224 xm1224 2.99137106960636e-14
Vx1224 xm1224 0 0
Gx1224_2 x1224 0 u2 0 -1.46395168088294e-08
Rx1225 x1225 0 1
Fxc1225_1224 x1225 0 Vx1224 -687.645107066235
Cx1225 x1225 xm1225 2.99137106960636e-14
Vx1225 xm1225 0 0
Gx1225_2 x1225 0 u2 0 1.00667921034054e-05
Rx1226 x1226 0 1
Fxc1226_1227 x1226 0 Vx1227 155.167635159053
Cx1226 x1226 xm1226 2.79263378446223e-13
Vx1226 xm1226 0 0
Gx1226_2 x1226 0 u2 0 -3.15550007305176e-05
Rx1227 x1227 0 1
Fxc1227_1226 x1227 0 Vx1226 -95.9036602768841
Cx1227 x1227 xm1227 2.79263378446224e-13
Vx1227 xm1227 0 0
Gx1227_2 x1227 0 u2 0 0.00302624007009638
Rx1228 x1228 0 1
Fxc1228_1229 x1228 0 Vx1229 264.458060116817
Cx1228 x1228 xm1228 1.23092401377661e-13
Vx1228 xm1228 0 0
Gx1228_2 x1228 0 u2 0 -4.24280577816601e-06
Rx1229 x1229 0 1
Fxc1229_1228 x1229 0 Vx1228 -285.273082614739
Cx1229 x1229 xm1229 1.23092401377661e-13
Vx1229 xm1229 0 0
Gx1229_2 x1229 0 u2 0 0.00121035828327304
Rx1230 x1230 0 1
Fxc1230_1231 x1230 0 Vx1231 6.48153364186914
Cx1230 x1230 xm1230 2.82424764335851e-12
Vx1230 xm1230 0 0
Gx1230_2 x1230 0 u2 0 -0.0105471309357489
Rx1231 x1231 0 1
Fxc1231_1230 x1231 0 Vx1230 -25.152394277784
Cx1231 x1231 xm1231 2.82424764335851e-12
Vx1231 xm1231 0 0
Gx1231_2 x1231 0 u2 0 0.265285595795369
Rx1232 x1232 0 1
Fxc1232_1233 x1232 0 Vx1233 533.915482396108
Cx1232 x1232 xm1232 1.22590423162195e-13
Vx1232 xm1232 0 0
Gx1232_2 x1232 0 u2 0 -2.09662497745596e-06
Rx1233 x1233 0 1
Fxc1233_1232 x1233 0 Vx1232 -153.095632912126
Cx1233 x1233 xm1233 1.22590423162195e-13
Vx1233 xm1233 0 0
Gx1233_2 x1233 0 u2 0 0.000320984127902992
Rx1234 x1234 0 1
Fxc1234_1235 x1234 0 Vx1235 392.986382267722
Cx1234 x1234 xm1234 4.09020191567389e-13
Vx1234 xm1234 0 0
Gx1234_2 x1234 0 u2 0 -0.000118221262876462
Rx1235 x1235 0 1
Fxc1235_1234 x1235 0 Vx1234 -18.5906279404846
Cx1235 x1235 xm1235 4.09020191567389e-13
Vx1235 xm1235 0 0
Gx1235_2 x1235 0 u2 0 0.00219780751279054
Rx1236 x1236 0 1
Fxc1236_1237 x1236 0 Vx1237 3655.3048430659
Cx1236 x1236 xm1236 9.93705359088137e-14
Vx1236 xm1236 0 0
Gx1236_2 x1236 0 u2 0 -1.64741623433466e-06
Rx1237 x1237 0 1
Fxc1237_1236 x1237 0 Vx1236 -33.3695789714479
Cx1237 x1237 xm1237 9.93705359088137e-14
Vx1237 xm1237 0 0
Gx1237_2 x1237 0 u2 0 5.49735861304759e-05
Rx1238 x1238 0 1
Fxc1238_1239 x1238 0 Vx1239 504.542610830624
Cx1238 x1238 xm1238 5.79622437737296e-14
Vx1238 xm1238 0 0
Gx1238_2 x1238 0 u2 0 -1.66428651606889e-07
Rx1239 x1239 0 1
Fxc1239_1238 x1239 0 Vx1238 -685.09336483455
Cx1239 x1239 xm1239 5.79622437737296e-14
Vx1239 xm1239 0 0
Gx1239_2 x1239 0 u2 0 0.000114019164934241
Rx1240 x1240 0 1
Fxc1240_1241 x1240 0 Vx1241 19935.8779799908
Cx1240 x1240 xm1240 3.54576514760153e-14
Vx1240 xm1240 0 0
Gx1240_2 x1240 0 u2 0 -6.80455767986286e-08
Rx1241 x1241 0 1
Fxc1241_1240 x1241 0 Vx1240 -47.1665785557395
Cx1241 x1241 xm1241 3.54576514760153e-14
Vx1241 xm1241 0 0
Gx1241_2 x1241 0 u2 0 3.20947704344312e-06
Rx1242 x1242 0 1
Fxc1242_1243 x1242 0 Vx1243 92.0492523309302
Cx1242 x1242 xm1242 1.2896763528379e-13
Vx1242 xm1242 0 0
Gx1242_2 x1242 0 u2 0 -1.21282294504326e-06
Rx1243 x1243 0 1
Fxc1243_1242 x1243 0 Vx1242 -782.055549819662
Cx1243 x1243 xm1243 1.2896763528379e-13
Vx1243 xm1243 0 0
Gx1243_2 x1243 0 u2 0 0.000948494915119711
Rx1244 x1244 0 1
Fxc1244_1245 x1244 0 Vx1245 469.912871689852
Cx1244 x1244 xm1244 9.26424551985641e-14
Vx1244 xm1244 0 0
Gx1244_2 x1244 0 u2 0 -6.81094118703232e-07
Rx1245 x1245 0 1
Fxc1245_1244 x1245 0 Vx1244 -307.781681490112
Cx1245 x1245 xm1245 9.26424551985641e-14
Vx1245 xm1245 0 0
Gx1245_2 x1245 0 u2 0 0.000209628293107506
Rx1246 x1246 0 1
Fxc1246_1247 x1246 0 Vx1247 5617.0715812471
Cx1246 x1246 xm1246 1.72944646712239e-14
Vx1246 xm1246 0 0
Gx1246_2 x1246 0 u2 0 -1.55980588421271e-08
Rx1247 x1247 0 1
Fxc1247_1246 x1247 0 Vx1246 -745.871639032922
Cx1247 x1247 xm1247 1.72944646712239e-14
Vx1247 xm1247 0 0
Gx1247_2 x1247 0 u2 0 1.16341497143093e-05
Rx1248 x1248 0 1
Fxc1248_1249 x1248 0 Vx1249 29.9082733827951
Cx1248 x1248 xm1248 3.11153675188471e-13
Vx1248 xm1248 0 0
Gx1248_2 x1248 0 u2 0 -4.03001523570316e-06
Rx1249 x1249 0 1
Fxc1249_1248 x1249 0 Vx1248 -482.764805045078
Cx1249 x1249 xm1249 3.11153675188471e-13
Vx1249 xm1249 0 0
Gx1249_2 x1249 0 u2 0 0.00194554951959293
Rx1250 x1250 0 1
Fxc1250_1251 x1250 0 Vx1251 89.7629700398008
Cx1250 x1250 xm1250 4.37725075845039e-13
Vx1250 xm1250 0 0
Gx1250_2 x1250 0 u2 0 -5.41771306322633e-05
Rx1251 x1251 0 1
Fxc1251_1250 x1251 0 Vx1250 -79.569779522322
Cx1251 x1251 xm1251 4.37725075845039e-13
Vx1251 xm1251 0 0
Gx1251_2 x1251 0 u2 0 0.00431086233956123
Rx1252 x1252 0 1
Fxc1252_1253 x1252 0 Vx1253 8.84393338199494
Cx1252 x1252 xm1252 2.89789505961041e-14
Vx1252 xm1252 0 0
Gx1252_2 x1252 0 u2 0 -2.71840711809331e-10
Rx1253 x1253 0 1
Fxc1253_1252 x1253 0 Vx1252 -172229.172750429
Cx1253 x1253 xm1253 2.89789505961041e-14
Vx1253 xm1253 0 0
Gx1253_2 x1253 0 u2 0 4.68189009148089e-05
Rx1254 x1254 0 1
Fxc1254_1255 x1254 0 Vx1255 59.898478011566
Cx1254 x1254 xm1254 3.08257267736937e-13
Vx1254 xm1254 0 0
Gx1254_2 x1254 0 u2 0 -1.07450037744446e-05
Rx1255 x1255 0 1
Fxc1255_1254 x1255 0 Vx1254 -231.419509563122
Cx1255 x1255 xm1255 3.08257267736937e-13
Vx1255 xm1255 0 0
Gx1255_2 x1255 0 u2 0 0.00248660350373587
Rx1256 x1256 0 1
Fxc1256_1257 x1256 0 Vx1257 2904.32747621958
Cx1256 x1256 xm1256 6.93829485175084e-14
Vx1256 xm1256 0 0
Gx1256_2 x1256 0 u2 0 -2.50043819806951e-07
Rx1257 x1257 0 1
Fxc1257_1256 x1257 0 Vx1256 -92.7711348607296
Cx1257 x1257 xm1257 6.93829485175084e-14
Vx1257 xm1257 0 0
Gx1257_2 x1257 0 u2 0 2.31968489284026e-05
Rx1258 x1258 0 1
Fxc1258_1259 x1258 0 Vx1259 78.8304304688954
Cx1258 x1258 xm1258 8.93653863244677e-14
Vx1258 xm1258 0 0
Gx1258_2 x1258 0 u2 0 -8.95592112107164e-08
Rx1259 x1259 0 1
Fxc1259_1258 x1259 0 Vx1258 -2161.33046187128
Cx1259 x1259 xm1259 8.93653863244677e-14
Vx1259 xm1259 0 0
Gx1259_2 x1259 0 u2 0 0.000193567051330885
Rx1260 x1260 0 1
Fxc1260_1261 x1260 0 Vx1261 947.937658111715
Cx1260 x1260 xm1260 7.05517351858277e-14
Vx1260 xm1260 0 0
Gx1260_2 x1260 0 u2 0 -2.6537122803651e-07
Rx1261 x1261 0 1
Fxc1261_1260 x1261 0 Vx1260 -277.354578049794
Cx1261 x1261 xm1261 7.05517351858277e-14
Vx1261 xm1261 0 0
Gx1261_2 x1261 0 u2 0 7.3601924978622e-05
Rx1262 x1262 0 1
Fxc1262_1263 x1262 0 Vx1263 2951.85320451397
Cx1262 x1262 xm1262 1.82509464382829e-14
Vx1262 xm1262 0 0
Gx1262_2 x1262 0 u2 0 -9.53240236698459e-09
Rx1263 x1263 0 1
Fxc1263_1262 x1263 0 Vx1262 -1398.31067098214
Cx1263 x1263 xm1263 1.82509464382829e-14
Vx1263 xm1263 0 0
Gx1263_2 x1263 0 u2 0 1.33292599498499e-05
Rx1264 x1264 0 1
Fxc1264_1265 x1264 0 Vx1265 1822.67872309301
Cx1264 x1264 xm1264 2.53969224170102e-14
Vx1264 xm1264 0 0
Gx1264_2 x1264 0 u2 0 -2.56468592779997e-08
Rx1265 x1265 0 1
Fxc1265_1264 x1265 0 Vx1264 -1131.14066462744
Cx1265 x1265 xm1265 2.53969224170102e-14
Vx1265 xm1265 0 0
Gx1265_2 x1265 0 u2 0 2.90102054493228e-05
Rx1266 x1266 0 1
Fxc1266_1267 x1266 0 Vx1267 6772.38611878903
Cx1266 x1266 xm1266 2.15604352286955e-14
Vx1266 xm1266 0 0
Gx1266_2 x1266 0 u2 0 -2.39543705459431e-08
Rx1267 x1267 0 1
Fxc1267_1266 x1267 0 Vx1266 -447.732368084428
Cx1267 x1267 xm1267 2.15604352286955e-14
Vx1267 xm1267 0 0
Gx1267_2 x1267 0 u2 0 1.0725147050507e-05
Rx1268 x1268 0 1
Fxc1268_1269 x1268 0 Vx1269 2.62148615304885
Cx1268 x1268 xm1268 6.88076389610427e-14
Vx1268 xm1268 0 0
Gx1268_2 x1268 0 u2 0 -7.49682497724048e-10
Rx1269 x1269 0 1
Fxc1269_1268 x1269 0 Vx1268 -115144.926755536
Cx1269 x1269 xm1269 6.88076389610427e-14
Vx1269 xm1269 0 0
Gx1269_2 x1269 0 u2 0 8.63221362903429e-05
Rx1270 x1270 0 1
Fxc1270_1271 x1270 0 Vx1271 657.979191374933
Cx1270 x1270 xm1270 3.36224705594798e-14
Vx1270 xm1270 0 0
Gx1270_2 x1270 0 u2 0 -1.9804683170983e-08
Rx1271 x1271 0 1
Fxc1271_1270 x1271 0 Vx1270 -1944.73484654513
Cx1271 x1271 xm1271 3.36224705594798e-14
Vx1271 xm1271 0 0
Gx1271_2 x1271 0 u2 0 3.85148574873965e-05
Rx1272 x1272 0 1
Fxc1272_1273 x1272 0 Vx1273 431.00516572359
Cx1272 x1272 xm1272 3.82271448805577e-14
Vx1272 xm1272 0 0
Gx1272_2 x1272 0 u2 0 -1.45185578368648e-08
Rx1273 x1273 0 1
Fxc1273_1272 x1273 0 Vx1272 -2342.78102221939
Cx1273 x1273 xm1273 3.82271448805577e-14
Vx1273 xm1273 0 0
Gx1273_2 x1273 0 u2 0 3.40138017702014e-05
Rx1274 x1274 0 1
Fxc1274_1275 x1274 0 Vx1275 30.3125416372388
Cx1274 x1274 xm1274 1.20061702453183e-13
Vx1274 xm1274 0 0
Gx1274_2 x1274 0 u2 0 -8.71978082219806e-08
Rx1275 x1275 0 1
Fxc1275_1274 x1275 0 Vx1274 -3448.41973580158
Cx1275 x1275 xm1275 1.20061702453183e-13
Vx1275 xm1275 0 0
Gx1275_2 x1275 0 u2 0 0.000300694642791319
Rx1276 x1276 0 1
Fxc1276_1277 x1276 0 Vx1277 2752.54685607216
Cx1276 x1276 xm1276 5.54932867986001e-14
Vx1276 xm1276 0 0
Gx1276_2 x1276 0 u2 0 -1.22446941227606e-07
Rx1277 x1277 0 1
Fxc1277_1276 x1277 0 Vx1276 -176.609190425089
Cx1277 x1277 xm1277 5.54932867986001e-14
Vx1277 xm1277 0 0
Gx1277_2 x1277 0 u2 0 2.16252551602359e-05
Rx1278 x1278 0 1
Fxc1278_1279 x1278 0 Vx1279 380.555191420678
Cx1278 x1278 xm1278 6.24009086699586e-14
Vx1278 xm1278 0 0
Gx1278_2 x1278 0 u2 0 -1.01377754934628e-07
Rx1279 x1279 0 1
Fxc1279_1278 x1279 0 Vx1278 -1028.24299254141
Cx1279 x1279 xm1279 6.24009086699586e-14
Vx1279 xm1279 0 0
Gx1279_2 x1279 0 u2 0 0.000104240966111111
Rx1280 x1280 0 1
Fxc1280_1281 x1280 0 Vx1281 50.3615745082337
Cx1280 x1280 xm1280 6.64567064981729e-14
Vx1280 xm1280 0 0
Gx1280_2 x1280 0 u2 0 -1.99629197074502e-08
Rx1281 x1281 0 1
Fxc1281_1280 x1281 0 Vx1280 -6893.29264876557
Cx1281 x1281 xm1281 6.64567064981729e-14
Vx1281 xm1281 0 0
Gx1281_2 x1281 0 u2 0 0.000137610247667264
Rx1282 x1282 0 1
Fxc1282_1283 x1282 0 Vx1283 78.2678260141868
Cx1282 x1282 xm1282 1.92779692469307e-13
Vx1282 xm1282 0 0
Gx1282_2 x1282 0 u2 0 -1.05095167548822e-06
Rx1283 x1283 0 1
Fxc1283_1282 x1283 0 Vx1282 -535.795986764311
Cx1283 x1283 xm1283 1.92779692469307e-13
Vx1283 xm1283 0 0
Gx1283_2 x1283 0 u2 0 0.000563095690009814
Rx1284 x1284 0 1
Fxc1284_1285 x1284 0 Vx1285 174.738554021833
Cx1284 x1284 xm1284 1.15282449142532e-12
Vx1284 xm1284 0 0
Gx1284_2 x1284 0 u2 0 -0.00035830080011358
Rx1285 x1285 0 1
Fxc1285_1284 x1285 0 Vx1284 -7.46531515671294
Cx1285 x1285 xm1285 1.15282449142532e-12
Vx1285 xm1285 0 0
Gx1285_2 x1285 0 u2 0 0.00267482839375028
Rx1286 x1286 0 1
Fxc1286_1287 x1286 0 Vx1287 1024.16634202391
Cx1286 x1286 xm1286 2.87628016359056e-14
Vx1286 xm1286 0 0
Gx1286_2 x1286 0 u2 0 -1.47602369459525e-08
Rx1287 x1287 0 1
Fxc1287_1286 x1287 0 Vx1286 -1845.34843575769
Cx1287 x1287 xm1287 2.87628016359056e-14
Vx1287 xm1287 0 0
Gx1287_2 x1287 0 u2 0 2.72377801596262e-05
Rx1288 x1288 0 1
Fxc1288_1289 x1288 0 Vx1289 18.4386393563261
Cx1288 x1288 xm1288 1.78666875824597e-13
Vx1288 xm1288 0 0
Gx1288_2 x1288 0 u2 0 -1.64995627098761e-07
Rx1289 x1289 0 1
Fxc1289_1288 x1289 0 Vx1288 -2717.03218370115
Cx1289 x1289 xm1289 1.78666875824597e-13
Vx1289 xm1289 0 0
Gx1289_2 x1289 0 u2 0 0.000448298428997288
Rx1290 x1290 0 1
Fxc1290_1291 x1290 0 Vx1291 957.050839521842
Cx1290 x1290 xm1290 1.04155247034917e-13
Vx1290 xm1290 0 0
Gx1290_2 x1290 0 u2 0 -4.63567202711241e-07
Rx1291 x1291 0 1
Fxc1291_1290 x1291 0 Vx1290 -152.860019763419
Cx1291 x1291 xm1291 1.04155247034917e-13
Vx1291 xm1291 0 0
Gx1291_2 x1291 0 u2 0 7.08608917681132e-05
Rx1292 x1292 0 1
Fxc1292_1293 x1292 0 Vx1293 6555.28728972687
Cx1292 x1292 xm1292 1.06235443062179e-14
Vx1292 xm1292 0 0
Gx1292_2 x1292 0 u2 0 -4.53210125618578e-09
Rx1293 x1293 0 1
Fxc1293_1292 x1293 0 Vx1292 -2203.62741654336
Cx1293 x1293 xm1293 1.06235443062179e-14
Vx1293 xm1293 0 0
Gx1293_2 x1293 0 u2 0 9.98706258268159e-06
Rx1294 x1294 0 1
Fxc1294_1295 x1294 0 Vx1295 504.724131461466
Cx1294 x1294 xm1294 5.41238890095385e-14
Vx1294 xm1294 0 0
Gx1294_2 x1294 0 u2 0 -2.47894475760694e-08
Rx1295 x1295 0 1
Fxc1295_1294 x1295 0 Vx1294 -1121.71262091002
Cx1295 x1295 xm1295 5.41238890095385e-14
Vx1295 xm1295 0 0
Gx1295_2 x1295 0 u2 0 2.78066362114643e-05
Rx1296 x1296 0 1
Fxc1296_1297 x1296 0 Vx1297 879.73452901079
Cx1296 x1296 xm1296 3.3864832840636e-14
Vx1296 xm1296 0 0
Gx1296_2 x1296 0 u2 0 -2.09736120679723e-08
Rx1297 x1297 0 1
Fxc1297_1296 x1297 0 Vx1296 -1661.46310520591
Cx1297 x1297 xm1297 3.3864832840636e-14
Vx1297 xm1297 0 0
Gx1297_2 x1297 0 u2 0 3.48468826338374e-05
Rx1298 x1298 0 1
Fxc1298_1299 x1298 0 Vx1299 24.2184135190404
Cx1298 x1298 xm1298 4.1684778621004e-13
Vx1298 xm1298 0 0
Gx1298_2 x1298 0 u2 0 -5.42987426355481e-06
Rx1299 x1299 0 1
Fxc1299_1298 x1299 0 Vx1298 -419.472146318784
Cx1299 x1299 xm1299 4.1684778621004e-13
Vx1299 xm1299 0 0
Gx1299_2 x1299 0 u2 0 0.00227768101157446
Rx1300 x1300 0 1
Fxc1300_1301 x1300 0 Vx1301 450.370392538576
Cx1300 x1300 xm1300 1.43290144219323e-14
Vx1300 xm1300 0 0
Gx1300_2 x1300 0 u2 0 -9.32132274181779e-10
Rx1301 x1301 0 1
Fxc1301_1300 x1301 0 Vx1300 -18561.04142872
Cx1301 x1301 xm1301 1.43290144219323e-14
Vx1301 xm1301 0 0
Gx1301_2 x1301 0 u2 0 1.7301345758135e-05
Rx1302 x1302 0 1
Fxc1302_1303 x1302 0 Vx1303 6062.70218589461
Cx1302 x1302 xm1302 1.59153780242877e-14
Vx1302 xm1302 0 0
Gx1302_2 x1302 0 u2 0 -2.08508137505182e-09
Rx1303 x1303 0 1
Fxc1303_1302 x1303 0 Vx1302 -1187.96000640292
Cx1303 x1303 xm1303 1.59153780242877e-14
Vx1303 xm1303 0 0
Gx1303_2 x1303 0 u2 0 2.47699328365717e-06
Rx1304 x1304 0 1
Fxc1304_1305 x1304 0 Vx1305 1220.43825025268
Cx1304 x1304 xm1304 1.1293667793922e-13
Vx1304 xm1304 0 0
Gx1304_2 x1304 0 u2 0 -3.57685591495425e-07
Rx1305 x1305 0 1
Fxc1305_1304 x1305 0 Vx1304 -116.154816172404
Cx1305 x1305 xm1305 1.1293667793922e-13
Vx1305 xm1305 0 0
Gx1305_2 x1305 0 u2 0 4.15469041276687e-05
Rx1306 x1306 0 1
Fxc1306_1307 x1306 0 Vx1307 817.776015036308
Cx1306 x1306 xm1306 1.00794993851598e-13
Vx1306 xm1306 0 0
Gx1306_2 x1306 0 u2 0 -3.84356722451948e-07
Rx1307 x1307 0 1
Fxc1307_1306 x1307 0 Vx1306 -214.414041963294
Cx1307 x1307 xm1307 1.00794993851598e-13
Vx1307 xm1307 0 0
Gx1307_2 x1307 0 u2 0 8.24114784166862e-05
Rx1308 x1308 0 1
Fxc1308_1309 x1308 0 Vx1309 197.197117286454
Cx1308 x1308 xm1308 3.93436377555167e-14
Vx1308 xm1308 0 0
Gx1308_2 x1308 0 u2 0 -6.13948923542168e-09
Rx1309 x1309 0 1
Fxc1309_1308 x1309 0 Vx1308 -5759.53272360174
Cx1309 x1309 xm1309 3.93436377555167e-14
Vx1309 xm1309 0 0
Gx1309_2 x1309 0 u2 0 3.53605891576118e-05
Rx1310 x1310 0 1
Fxc1310_1311 x1310 0 Vx1311 2883.56987994648
Cx1310 x1310 xm1310 4.27323643580748e-14
Vx1310 xm1310 0 0
Gx1310_2 x1310 0 u2 0 -1.37905519088704e-08
Rx1311 x1311 0 1
Fxc1311_1310 x1311 0 Vx1310 -354.894212503292
Cx1311 x1311 xm1311 4.27323643580748e-14
Vx1311 xm1311 0 0
Gx1311_2 x1311 0 u2 0 4.89418705968432e-06
Rx1312 x1312 0 1
Cx1312 x1312 0 1.40144076963712e-10
Gx1312_2 x1312 0 u2 0 -38.1873028477036
Rx1313 x1313 0 1
Fxc1313_1314 x1313 0 Vx1314 44.7040859600632
Cx1313 x1313 xm1313 1.39431711841145e-12
Vx1313 xm1313 0 0
Gx1313_2 x1313 0 u2 0 -0.000606850354415158
Rx1314 x1314 0 1
Fxc1314_1313 x1314 0 Vx1313 -24.8558273951751
Cx1314 x1314 xm1314 1.39431711841145e-12
Vx1314 xm1314 0 0
Gx1314_2 x1314 0 u2 0 0.015083767664044
Rx1315 x1315 0 1
Fxc1315_1316 x1315 0 Vx1316 14660.6684346308
Cx1315 x1315 xm1315 4.46055376469595e-14
Vx1315 xm1315 0 0
Gx1315_2 x1315 0 u2 0 -3.92432706306805e-08
Rx1316 x1316 0 1
Fxc1316_1315 x1316 0 Vx1315 -70.5798265469312
Cx1316 x1316 xm1316 4.46055376469595e-14
Vx1316 xm1316 0 0
Gx1316_2 x1316 0 u2 0 2.76978323424771e-06
Rx1317 x1317 0 1
Fxc1317_1318 x1317 0 Vx1318 186.685134523892
Cx1317 x1317 xm1317 1.38311295911203e-13
Vx1317 xm1317 0 0
Gx1317_2 x1317 0 u2 0 -9.44568304252493e-07
Rx1318 x1318 0 1
Fxc1318_1317 x1318 0 Vx1317 -557.098521823304
Cx1318 x1318 xm1318 1.38311295911203e-13
Vx1318 xm1318 0 0
Gx1318_2 x1318 0 u2 0 0.000526217606060208
Rx1319 x1319 0 1
Fxc1319_1320 x1319 0 Vx1320 8.10107632863315
Cx1319 x1319 xm1319 2.19578957008743e-13
Vx1319 xm1319 0 0
Gx1319_2 x1319 0 u2 0 -2.39461227263102e-07
Rx1320 x1320 0 1
Fxc1320_1319 x1320 0 Vx1319 -5104.32447619449
Cx1320 x1320 xm1320 2.19578957008743e-13
Vx1320 xm1320 0 0
Gx1320_2 x1320 0 u2 0 0.00122228780341862
Rx1321 x1321 0 1
Fxc1321_1322 x1321 0 Vx1322 977.765602899993
Cx1321 x1321 xm1321 4.73505553997717e-14
Vx1321 xm1321 0 0
Gx1321_2 x1321 0 u2 0 -1.90480814329219e-08
Rx1322 x1322 0 1
Fxc1322_1321 x1322 0 Vx1321 -870.685647413662
Cx1322 x1322 xm1322 4.73505553997717e-14
Vx1322 xm1322 0 0
Gx1322_2 x1322 0 u2 0 1.65848911144118e-05
Rx1323 x1323 0 1
Fxc1323_1324 x1323 0 Vx1324 212.19164058068
Cx1323 x1323 xm1323 1.22056182242707e-13
Vx1323 xm1323 0 0
Gx1323_2 x1323 0 u2 0 -2.03824609815998e-07
Rx1324 x1324 0 1
Fxc1324_1323 x1324 0 Vx1323 -611.616455380204
Cx1324 x1324 xm1324 1.22056182242707e-13
Vx1324 xm1324 0 0
Gx1324_2 x1324 0 u2 0 0.000124662485374914
Rx1325 x1325 0 1
Fxc1325_1326 x1325 0 Vx1326 1867.81786279149
Cx1325 x1325 xm1325 4.2540439057887e-14
Vx1325 xm1325 0 0
Gx1325_2 x1325 0 u2 0 -4.2488561497154e-08
Rx1326 x1326 0 1
Fxc1326_1325 x1326 0 Vx1325 -579.865590923381
Cx1326 x1326 xm1326 4.2540439057887e-14
Vx1326 xm1326 0 0
Gx1326_2 x1326 0 u2 0 2.46376548200316e-05
Rx1327 x1327 0 1
Fxc1327_1328 x1327 0 Vx1328 0.552506355563814
Cx1327 x1327 xm1327 8.16769439323924e-11
Vx1327 xm1327 0 0
Gx1327_2 x1327 0 u2 0 -16.8453383263521
Rx1328 x1328 0 1
Fxc1328_1327 x1328 0 Vx1327 -1.23156497795124
Cx1328 x1328 xm1328 8.16769439323924e-11
Vx1328 xm1328 0 0
Gx1328_2 x1328 0 u2 0 20.7461287244751
Rx1329 x1329 0 1
Fxc1329_1330 x1329 0 Vx1330 0.201922100496264
Cx1329 x1329 xm1329 3.055355601781e-12
Vx1329 xm1329 0 0
Gx1329_2 x1329 0 u2 0 -6.19838416591743e-05
Rx1330 x1330 0 1
Fxc1330_1329 x1330 0 Vx1329 -1303.75549727767
Cx1330 x1330 xm1330 3.055355601781e-12
Vx1330 xm1330 0 0
Gx1330_2 x1330 0 u2 0 0.0808117743055375
Rx1331 x1331 0 1
Fxc1331_1332 x1331 0 Vx1332 10.2931396678079
Cx1331 x1331 xm1331 2.22336076590458e-13
Vx1331 xm1331 0 0
Gx1331_2 x1331 0 u2 0 -9.79281880341221e-08
Rx1332 x1332 0 1
Fxc1332_1331 x1332 0 Vx1331 -4847.45705959316
Cx1332 x1332 xm1332 2.22336076590458e-13
Vx1332 xm1332 0 0
Gx1332_2 x1332 0 u2 0 0.000474702686419172
Rx1333 x1333 0 1
Fxc1333_1334 x1333 0 Vx1334 49.2732062416815
Cx1333 x1333 xm1333 7.0682437690172e-13
Vx1333 xm1333 0 0
Gx1333_2 x1333 0 u2 0 -4.87201457186929e-05
Rx1334 x1334 0 1
Fxc1334_1333 x1334 0 Vx1333 -90.7364887247144
Cx1334 x1334 xm1334 7.0682437690172e-13
Vx1334 xm1334 0 0
Gx1334_2 x1334 0 u2 0 0.00442069495267062
Rx1335 x1335 0 1
Fxc1335_1336 x1335 0 Vx1336 195.955468404239
Cx1335 x1335 xm1335 5.1045195384584e-14
Vx1335 xm1335 0 0
Gx1335_2 x1335 0 u2 0 -1.20068446604254e-08
Rx1336 x1336 0 1
Fxc1336_1335 x1336 0 Vx1335 -4097.88927995572
Cx1336 x1336 xm1336 5.1045195384584e-14
Vx1336 xm1336 0 0
Gx1336_2 x1336 0 u2 0 4.92027200200507e-05
Rx1337 x1337 0 1
Fxc1337_1338 x1337 0 Vx1338 857.728958787232
Cx1337 x1337 xm1337 2.41223264060163e-13
Vx1337 xm1337 0 0
Gx1337_2 x1337 0 u2 0 -2.0439071681426e-06
Rx1338 x1338 0 1
Fxc1338_1337 x1338 0 Vx1337 -43.0072668806513
Cx1338 x1338 xm1338 2.41223264060163e-13
Vx1338 xm1338 0 0
Gx1338_2 x1338 0 u2 0 8.7902861059585e-05
Rx1339 x1339 0 1
Fxc1339_1340 x1339 0 Vx1340 2801.70460222655
Cx1339 x1339 xm1339 9.93476076097149e-14
Vx1339 xm1339 0 0
Gx1339_2 x1339 0 u2 0 -1.78669550173755e-07
Rx1340 x1340 0 1
Fxc1340_1339 x1340 0 Vx1339 -78.8169791687942
Cx1340 x1340 xm1340 9.93476076097149e-14
Vx1340 xm1340 0 0
Gx1340_2 x1340 0 u2 0 1.40821942141427e-05
Rx1341 x1341 0 1
Fxc1341_1342 x1341 0 Vx1342 1997.19587059298
Cx1341 x1341 xm1341 1.96255535649835e-14
Vx1341 xm1341 0 0
Gx1341_2 x1341 0 u2 0 -7.71567535262718e-09
Rx1342 x1342 0 1
Fxc1342_1341 x1342 0 Vx1341 -2910.21753683064
Cx1342 x1342 xm1342 1.96255535649835e-14
Vx1342 xm1342 0 0
Gx1342_2 x1342 0 u2 0 2.24542937197076e-05
Rx1343 x1343 0 1
Fxc1343_1344 x1343 0 Vx1344 217.922987869194
Cx1343 x1343 xm1343 2.15369618623669e-13
Vx1343 xm1343 0 0
Gx1343_2 x1343 0 u2 0 -1.03655083220309e-06
Rx1344 x1344 0 1
Fxc1344_1343 x1344 0 Vx1343 -227.275981907037
Cx1344 x1344 xm1344 2.15369618623669e-13
Vx1344 xm1344 0 0
Gx1344_2 x1344 0 u2 0 0.000235583108185514
Rx1345 x1345 0 1
Fxc1345_1346 x1345 0 Vx1346 4017.04261481846
Cx1345 x1345 xm1345 1.21891798583539e-14
Vx1345 xm1345 0 0
Gx1345_2 x1345 0 u2 0 -8.6557728772054e-10
Rx1346 x1346 0 1
Fxc1346_1345 x1346 0 Vx1345 -3551.61707126844
Cx1346 x1346 xm1346 1.21891798583539e-14
Vx1346 xm1346 0 0
Gx1346_2 x1346 0 u2 0 3.0741990715705e-06
Rx1347 x1347 0 1
Fxc1347_1348 x1347 0 Vx1348 1324.11108100025
Cx1347 x1347 xm1347 2.69942236556942e-14
Vx1347 xm1347 0 0
Gx1347_2 x1347 0 u2 0 -9.67759747335958e-09
Rx1348 x1348 0 1
Fxc1348_1347 x1348 0 Vx1347 -2497.00825751769
Cx1348 x1348 xm1348 2.69942236556942e-14
Vx1348 xm1348 0 0
Gx1348_2 x1348 0 u2 0 2.41650408039113e-05
Rx1349 x1349 0 1
Fxc1349_1350 x1349 0 Vx1350 53.7733401901532
Cx1349 x1349 xm1349 7.7544284673081e-14
Vx1349 xm1349 0 0
Gx1349_2 x1349 0 u2 0 -6.54652583565449e-09
Rx1350 x1350 0 1
Fxc1350_1349 x1350 0 Vx1349 -7225.93697971421
Cx1350 x1350 xm1350 7.7544284673081e-14
Vx1350 xm1350 0 0
Gx1350_2 x1350 0 u2 0 4.73047831245103e-05
Rx1351 x1351 0 1
Fxc1351_1352 x1351 0 Vx1352 1274.87815290969
Cx1351 x1351 xm1351 1.03543939234814e-13
Vx1351 xm1351 0 0
Gx1351_2 x1351 0 u2 0 -1.56624323692179e-07
Rx1352 x1352 0 1
Fxc1352_1351 x1352 0 Vx1351 -173.973949638349
Cx1352 x1352 xm1352 1.03543939234814e-13
Vx1352 xm1352 0 0
Gx1352_2 x1352 0 u2 0 2.72485522021635e-05
Rx1353 x1353 0 1
Fxc1353_1354 x1353 0 Vx1354 3363.77878007121
Cx1353 x1353 xm1353 9.1674395278034e-14
Vx1353 xm1353 0 0
Gx1353_2 x1353 0 u2 0 -2.4367985568473e-07
Rx1354 x1354 0 1
Fxc1354_1353 x1354 0 Vx1353 -87.8235470628794
Cx1354 x1354 xm1354 9.1674395278034e-14
Vx1354 xm1354 0 0
Gx1354_2 x1354 0 u2 0 2.14008292740036e-05
Rx1355 x1355 0 1
Fxc1355_1356 x1355 0 Vx1356 359.594376381447
Cx1355 x1355 xm1355 1.90368710342961e-13
Vx1355 xm1355 0 0
Gx1355_2 x1355 0 u2 0 -8.26238355222181e-07
Rx1356 x1356 0 1
Fxc1356_1355 x1356 0 Vx1355 -196.738101631267
Cx1356 x1356 xm1356 1.90368710342961e-13
Vx1356 xm1356 0 0
Gx1356_2 x1356 0 u2 0 0.000162552565501352
Rx1357 x1357 0 1
Fxc1357_1358 x1357 0 Vx1358 889.86346713563
Cx1357 x1357 xm1357 3.43839976006569e-14
Vx1357 xm1357 0 0
Gx1357_2 x1357 0 u2 0 -9.79532500324516e-09
Rx1358 x1358 0 1
Fxc1358_1357 x1358 0 Vx1357 -2455.27629096701
Cx1358 x1358 xm1358 3.43839976006569e-14
Vx1358 xm1358 0 0
Gx1358_2 x1358 0 u2 0 2.40502292427842e-05
Rx1359 x1359 0 1
Fxc1359_1360 x1359 0 Vx1360 1687.12643990479
Cx1359 x1359 xm1359 1.10377999804161e-13
Vx1359 xm1359 0 0
Gx1359_2 x1359 0 u2 0 -1.24136362537118e-07
Rx1360 x1360 0 1
Fxc1360_1359 x1360 0 Vx1359 -127.725641914451
Cx1360 x1360 xm1360 1.10377999804161e-13
Vx1360 xm1360 0 0
Gx1360_2 x1360 0 u2 0 1.58553965899784e-05
Rx1361 x1361 0 1
Fxc1361_1362 x1361 0 Vx1362 1527.0860283956
Cx1361 x1361 xm1361 5.39843163452879e-14
Vx1361 xm1361 0 0
Gx1361_2 x1361 0 u2 0 -1.36080110482694e-08
Rx1362 x1362 0 1
Fxc1362_1361 x1362 0 Vx1361 -605.79619670411
Cx1362 x1362 xm1362 5.39843163452879e-14
Vx1362 xm1362 0 0
Gx1362_2 x1362 0 u2 0 8.24368133774913e-06
Rx1363 x1363 0 1
Fxc1363_1364 x1363 0 Vx1364 1043.78587254419
Cx1363 x1363 xm1363 1.66115615183985e-13
Vx1363 xm1363 0 0
Gx1363_2 x1363 0 u2 0 -4.31593480092347e-07
Rx1364 x1364 0 1
Fxc1364_1363 x1364 0 Vx1363 -95.0061762005637
Cx1364 x1364 xm1364 1.66115615183985e-13
Vx1364 xm1364 0 0
Gx1364_2 x1364 0 u2 0 4.1004046216668e-05
Rx1365 x1365 0 1
Fxc1365_1366 x1365 0 Vx1366 807.025070835754
Cx1365 x1365 xm1365 1.72753550245707e-13
Vx1365 xm1365 0 0
Gx1365_2 x1365 0 u2 0 -1.83743639135277e-06
Rx1366 x1366 0 1
Fxc1366_1365 x1366 0 Vx1365 -116.129570152787
Cx1366 x1366 xm1366 1.72753550245707e-13
Vx1366 xm1366 0 0
Gx1366_2 x1366 0 u2 0 0.000213380698310885
Rx1367 x1367 0 1
Fxc1367_1368 x1367 0 Vx1368 2893.32534377954
Cx1367 x1367 xm1367 7.89077374985022e-14
Vx1367 xm1367 0 0
Gx1367_2 x1367 0 u2 0 -2.97381838151889e-07
Rx1368 x1368 0 1
Fxc1368_1367 x1368 0 Vx1367 -155.150890802148
Cx1368 x1368 xm1368 7.89077374985021e-14
Vx1368 xm1368 0 0
Gx1368_2 x1368 0 u2 0 4.61390570976457e-05
Rx1369 x1369 0 1
Fxc1369_1370 x1369 0 Vx1370 37.5552030174587
Cx1369 x1369 xm1369 4.41676639181862e-13
Vx1369 xm1369 0 0
Gx1369_2 x1369 0 u2 0 -6.32061312527846e-06
Rx1370 x1370 0 1
Fxc1370_1369 x1370 0 Vx1369 -393.031883990262
Cx1370 x1370 xm1370 4.41676639181861e-13
Vx1370 xm1370 0 0
Gx1370_2 x1370 0 u2 0 0.00248420248460177
Rx1371 x1371 0 1
Fxc1371_1372 x1371 0 Vx1372 59.737267967888
Cx1371 x1371 xm1371 7.69508360165092e-13
Vx1371 xm1371 0 0
Gx1371_2 x1371 0 u2 0 -0.000284043284747505
Rx1372 x1372 0 1
Fxc1372_1371 x1372 0 Vx1371 -84.505006831606
Cx1372 x1372 xm1372 7.69508360165092e-13
Vx1372 xm1372 0 0
Gx1372_2 x1372 0 u2 0 0.0240030797180597
Rx1373 x1373 0 1
Fxc1373_1374 x1373 0 Vx1374 370.312705118759
Cx1373 x1373 xm1373 6.84174064919173e-13
Vx1373 xm1373 0 0
Gx1373_2 x1373 0 u2 0 -0.000445635151098327
Rx1374 x1374 0 1
Fxc1374_1373 x1374 0 Vx1373 -17.0599744999131
Cx1374 x1374 xm1374 6.84174064919173e-13
Vx1374 xm1374 0 0
Gx1374_2 x1374 0 u2 0 0.00760252431400239
Rx1375 x1375 0 1
Fxc1375_1376 x1375 0 Vx1376 540.998729506229
Cx1375 x1375 xm1375 3.41606667996328e-13
Vx1375 xm1375 0 0
Gx1375_2 x1375 0 u2 0 -2.21247183673026e-05
Rx1376 x1376 0 1
Fxc1376_1375 x1376 0 Vx1375 -46.7565970958917
Cx1376 x1376 xm1376 3.41606667996328e-13
Vx1376 xm1376 0 0
Gx1376_2 x1376 0 u2 0 0.00103447654256004
Rx1377 x1377 0 1
Fxc1377_1378 x1377 0 Vx1378 13.3875128016389
Cx1377 x1377 xm1377 1.07548830475537e-12
Vx1377 xm1377 0 0
Gx1377_2 x1377 0 u2 0 -3.90830105401504e-05
Rx1378 x1378 0 1
Fxc1378_1377 x1378 0 Vx1377 -204.611544257901
Cx1378 x1378 xm1378 1.07548830475537e-12
Vx1378 xm1378 0 0
Gx1378_2 x1378 0 u2 0 0.007996835140868
Rx1379 x1379 0 1
Fxc1379_1380 x1379 0 Vx1380 125.338908246659
Cx1379 x1379 xm1379 1.99049200010659e-13
Vx1379 xm1379 0 0
Gx1379_2 x1379 0 u2 0 -2.91820460125426e-07
Rx1380 x1380 0 1
Fxc1380_1379 x1380 0 Vx1379 -640.319514594647
Cx1380 x1380 xm1380 1.99049200010659e-13
Vx1380 xm1380 0 0
Gx1380_2 x1380 0 u2 0 0.000186858335376299
Rx1381 x1381 0 1
Fxc1381_1382 x1381 0 Vx1382 173.623366801763
Cx1381 x1381 xm1381 1.88237358199619e-13
Vx1381 xm1381 0 0
Gx1381_2 x1381 0 u2 0 -3.44112264609288e-07
Rx1382 x1382 0 1
Fxc1382_1381 x1382 0 Vx1381 -501.052685383336
Cx1382 x1382 xm1382 1.88237358199619e-13
Vx1382 xm1382 0 0
Gx1382_2 x1382 0 u2 0 0.000172418374255825
Rx1383 x1383 0 1
Fxc1383_1384 x1383 0 Vx1384 2602.59039055091
Cx1383 x1383 xm1383 1.57459489839352e-14
Vx1383 xm1383 0 0
Gx1383_2 x1383 0 u2 0 -2.0028745720622e-09
Rx1384 x1384 0 1
Fxc1384_1383 x1384 0 Vx1383 -4686.14721594799
Cx1384 x1384 xm1384 1.57459489839352e-14
Vx1384 xm1384 0 0
Gx1384_2 x1384 0 u2 0 9.38576509976233e-06
Rx1385 x1385 0 1
Fxc1385_1386 x1385 0 Vx1386 163036.839174037
Cx1385 x1385 xm1385 2.49001986220754e-14
Vx1385 xm1385 0 0
Gx1385_2 x1385 0 u2 0 -6.80351234202629e-09
Rx1386 x1386 0 1
Fxc1386_1385 x1386 0 Vx1385 -33.5687865766965
Cx1386 x1386 xm1386 2.49001986220754e-14
Vx1386 xm1386 0 0
Gx1386_2 x1386 0 u2 0 2.28385653781401e-07
Rx1387 x1387 0 1
Fxc1387_1388 x1387 0 Vx1388 101.538204423076
Cx1387 x1387 xm1387 1.20010327111104e-13
Vx1387 xm1387 0 0
Gx1387_2 x1387 0 u2 0 -3.24314618662399e-08
Rx1388 x1388 0 1
Fxc1388_1387 x1388 0 Vx1387 -2266.51264613607
Cx1388 x1388 xm1388 1.20010327111104e-13
Vx1388 xm1388 0 0
Gx1388_2 x1388 0 u2 0 7.35063184525124e-05
Rx1389 x1389 0 1
Fxc1389_1390 x1389 0 Vx1390 154.257543094607
Cx1389 x1389 xm1389 9.19589919698257e-13
Vx1389 xm1389 0 0
Gx1389_2 x1389 0 u2 0 -0.000154447735476183
Rx1390 x1390 0 1
Fxc1390_1389 x1390 0 Vx1389 -27.3399550494882
Cx1390 x1390 xm1390 9.19589919698257e-13
Vx1390 xm1390 0 0
Gx1390_2 x1390 0 u2 0 0.00422259414541408
Rx1391 x1391 0 1
Fxc1391_1392 x1391 0 Vx1392 135.434326759648
Cx1391 x1391 xm1391 1.35062615998325e-12
Vx1391 xm1391 0 0
Gx1391_2 x1391 0 u2 0 -0.000552561282987393
Rx1392 x1392 0 1
Fxc1392_1391 x1392 0 Vx1391 -14.4794141662475
Cx1392 x1392 xm1392 1.35062615998325e-12
Vx1392 xm1392 0 0
Gx1392_2 x1392 0 u2 0 0.00800076366860755
Rx1393 x1393 0 1
Fxc1393_1394 x1393 0 Vx1394 269197.10432815
Cx1393 x1393 xm1393 5.61403593569498e-16
Vx1393 xm1393 0 0
Gx1393_2 x1393 0 u2 0 -2.77517952406999e-10
Rx1394 x1394 0 1
Fxc1394_1393 x1394 0 Vx1393 -41235.6969749405
Cx1394 x1394 xm1394 5.61403593569498e-16
Vx1394 xm1394 0 0
Gx1394_2 x1394 0 u2 0 1.1443646190561e-05
Rx1395 x1395 0 1
Fxc1395_1396 x1395 0 Vx1396 141.682512324292
Cx1395 x1395 xm1395 1.34555540326277e-13
Vx1395 xm1395 0 0
Gx1395_2 x1395 0 u2 0 -8.43535856478129e-08
Rx1396 x1396 0 1
Fxc1396_1395 x1396 0 Vx1395 -1402.39299669797
Cx1396 x1396 xm1396 1.34555540326277e-13
Vx1396 xm1396 0 0
Gx1396_2 x1396 0 u2 0 0.000118296877758855
Rx1397 x1397 0 1
Fxc1397_1398 x1397 0 Vx1398 288.433733376754
Cx1397 x1397 xm1397 4.98865404960471e-13
Vx1397 xm1397 0 0
Gx1397_2 x1397 0 u2 0 -5.47540874929269e-06
Rx1398 x1398 0 1
Fxc1398_1397 x1398 0 Vx1397 -61.0431519566742
Cx1398 x1398 xm1398 4.98865404960471e-13
Vx1398 xm1398 0 0
Gx1398_2 x1398 0 u2 0 0.000334236208307977
Rx1399 x1399 0 1
Fxc1399_1400 x1399 0 Vx1400 79.7504425406474
Cx1399 x1399 xm1399 1.15714797739341e-12
Vx1399 xm1399 0 0
Gx1399_2 x1399 0 u2 0 -9.58574254610008e-05
Rx1400 x1400 0 1
Fxc1400_1399 x1400 0 Vx1399 -36.459645858532
Cx1400 x1400 xm1400 1.15714797739341e-12
Vx1400 xm1400 0 0
Gx1400_2 x1400 0 u2 0 0.00349492778521872
Rx1401 x1401 0 1
Fxc1401_1402 x1401 0 Vx1402 117.485744806806
Cx1401 x1401 xm1401 5.42048534221595e-13
Vx1401 xm1401 0 0
Gx1401_2 x1401 0 u2 0 -9.37143068718006e-06
Rx1402 x1402 0 1
Fxc1402_1401 x1402 0 Vx1401 -118.88643937028
Cx1402 x1402 xm1402 5.42048534221595e-13
Vx1402 xm1402 0 0
Gx1402_2 x1402 0 u2 0 0.00111413602620421
Rx1403 x1403 0 1
Fxc1403_1404 x1403 0 Vx1404 357.903216675792
Cx1403 x1403 xm1403 9.340099268043e-14
Vx1403 xm1403 0 0
Gx1403_2 x1403 0 u2 0 -5.45796154519508e-08
Rx1404 x1404 0 1
Fxc1404_1403 x1404 0 Vx1403 -1217.42886072467
Cx1404 x1404 xm1404 9.340099268043e-14
Vx1404 xm1404 0 0
Gx1404_2 x1404 0 u2 0 6.64467990584592e-05
Rx1405 x1405 0 1
Fxc1405_1406 x1405 0 Vx1406 422.431360853424
Cx1405 x1405 xm1405 2.02797650128333e-13
Vx1405 xm1405 0 0
Gx1405_2 x1405 0 u2 0 -4.40967383724686e-07
Rx1406 x1406 0 1
Fxc1406_1405 x1406 0 Vx1405 -242.844731438414
Cx1406 x1406 xm1406 2.02797650128333e-13
Vx1406 xm1406 0 0
Gx1406_2 x1406 0 u2 0 0.000107086605873722
Rx1407 x1407 0 1
Fxc1407_1408 x1407 0 Vx1408 69.4618475080829
Cx1407 x1407 xm1407 7.01742537232251e-13
Vx1407 xm1407 0 0
Gx1407_2 x1407 0 u2 0 -2.08408553199352e-05
Rx1408 x1408 0 1
Fxc1408_1407 x1408 0 Vx1407 -121.632654414284
Cx1408 x1408 xm1408 7.01742537232251e-13
Vx1408 xm1408 0 0
Gx1408_2 x1408 0 u2 0 0.00253492855282776
Rx1409 x1409 0 1
Fxc1409_1410 x1409 0 Vx1410 23.7338070751244
Cx1409 x1409 xm1409 6.4028082506253e-14
Vx1409 xm1409 0 0
Gx1409_2 x1409 0 u2 0 -1.55116426613005e-09
Rx1410 x1410 0 1
Fxc1410_1409 x1410 0 Vx1409 -38217.7287161464
Cx1410 x1410 xm1410 6.4028082506253e-14
Vx1410 xm1410 0 0
Gx1410_2 x1410 0 u2 0 5.92819751171385e-05
Rx1411 x1411 0 1
Fxc1411_1412 x1411 0 Vx1412 2169.50137004576
Cx1411 x1411 xm1411 3.68280434719191e-14
Vx1411 xm1411 0 0
Gx1411_2 x1411 0 u2 0 -2.02574681156965e-08
Rx1412 x1412 0 1
Fxc1412_1411 x1412 0 Vx1411 -1350.77467089874
Cx1412 x1412 xm1412 3.68280434719191e-14
Vx1412 xm1412 0 0
Gx1412_2 x1412 0 u2 0 2.73632748272217e-05
Rx1413 x1413 0 1
Fxc1413_1414 x1413 0 Vx1414 345.971584700494
Cx1413 x1413 xm1413 2.43463431944243e-13
Vx1413 xm1413 0 0
Gx1413_2 x1413 0 u2 0 -9.08346654293834e-07
Rx1414 x1414 0 1
Fxc1414_1413 x1414 0 Vx1413 -187.160837238373
Cx1414 x1414 xm1414 2.43463431944243e-13
Vx1414 xm1414 0 0
Gx1414_2 x1414 0 u2 0 0.000170006920320308
Rx1415 x1415 0 1
Fxc1415_1416 x1415 0 Vx1416 465.165456832328
Cx1415 x1415 xm1415 1.88338702913179e-13
Vx1415 xm1415 0 0
Gx1415_2 x1415 0 u2 0 -3.39186843018247e-07
Rx1416 x1416 0 1
Fxc1416_1415 x1416 0 Vx1415 -265.485675590252
Cx1416 x1416 xm1416 1.88338702913179e-13
Vx1416 xm1416 0 0
Gx1416_2 x1416 0 u2 0 9.00492481700238e-05
Rx1417 x1417 0 1
Fxc1417_1418 x1417 0 Vx1418 3959.71485741082
Cx1417 x1417 xm1417 4.99523803066435e-15
Vx1417 xm1417 0 0
Gx1417_2 x1417 0 u2 0 -7.26884916078383e-10
Rx1418 x1418 0 1
Fxc1418_1417 x1418 0 Vx1417 -45747.4860003254
Cx1418 x1418 xm1418 4.99523803066435e-15
Vx1418 xm1418 0 0
Gx1418_2 x1418 0 u2 0 3.32531575221435e-05
Rx1419 x1419 0 1
Fxc1419_1420 x1419 0 Vx1420 2.07826308785367
Cx1419 x1419 xm1419 7.43266824125504e-12
Vx1419 xm1419 0 0
Gx1419_2 x1419 0 u2 0 -0.00570764124292289
Rx1420 x1420 0 1
Fxc1420_1419 x1420 0 Vx1419 -51.5730176444532
Cx1420 x1420 xm1420 7.43266824125504e-12
Vx1420 xm1420 0 0
Gx1420_2 x1420 0 u2 0 0.294360282529471
Rx1421 x1421 0 1
Fxc1421_1422 x1421 0 Vx1422 31.8197370394212
Cx1421 x1421 xm1421 1.3706119903344e-12
Vx1421 xm1421 0 0
Gx1421_2 x1421 0 u2 0 -2.71690068954319e-05
Rx1422 x1422 0 1
Fxc1422_1421 x1422 0 Vx1421 -80.9999104186377
Cx1422 x1422 xm1422 1.3706119903344e-12
Vx1422 xm1422 0 0
Gx1422_2 x1422 0 u2 0 0.00220068712469333
Rx1423 x1423 0 1
Fxc1423_1424 x1423 0 Vx1424 2323.641248737
Cx1423 x1423 xm1423 1.32600732830319e-13
Vx1423 xm1423 0 0
Gx1423_2 x1423 0 u2 0 -1.25308170414251e-07
Rx1424 x1424 0 1
Fxc1424_1423 x1424 0 Vx1423 -115.993822312128
Cx1424 x1424 xm1424 1.32600732830319e-13
Vx1424 xm1424 0 0
Gx1424_2 x1424 0 u2 0 1.45349736532885e-05
Rx1425 x1425 0 1
Fxc1425_1426 x1425 0 Vx1426 896.240171386843
Cx1425 x1425 xm1425 6.7800124285245e-14
Vx1425 xm1425 0 0
Gx1425_2 x1425 0 u2 0 -1.7576663013938e-08
Rx1426 x1426 0 1
Fxc1426_1425 x1426 0 Vx1425 -1185.89112631769
Cx1426 x1426 xm1426 6.7800124285245e-14
Vx1426 xm1426 0 0
Gx1426_2 x1426 0 u2 0 2.08440086985055e-05
Rx1427 x1427 0 1
Fxc1427_1428 x1427 0 Vx1428 28.8085698038238
Cx1427 x1427 xm1427 1.115641621969e-13
Vx1427 xm1427 0 0
Gx1427_2 x1427 0 u2 0 -5.32601495290164e-09
Rx1428 x1428 0 1
Fxc1428_1427 x1428 0 Vx1427 -13924.6729789031
Cx1428 x1428 xm1428 1.115641621969e-13
Vx1428 xm1428 0 0
Gx1428_2 x1428 0 u2 0 7.41630164999036e-05
Rx1429 x1429 0 1
Fxc1429_1430 x1429 0 Vx1430 121.246729575124
Cx1429 x1429 xm1429 2.72702074238325e-13
Vx1429 xm1429 0 0
Gx1429_2 x1429 0 u2 0 -2.10375086357476e-07
Rx1430 x1430 0 1
Fxc1430_1429 x1430 0 Vx1429 -579.804116230625
Cx1430 x1430 xm1430 2.72702074238325e-13
Vx1430 xm1430 0 0
Gx1430_2 x1430 0 u2 0 0.000121976341022438
Rx1431 x1431 0 1
Fxc1431_1432 x1431 0 Vx1432 33.5755216439265
Cx1431 x1431 xm1431 1.01079656034734e-12
Vx1431 xm1431 0 0
Gx1431_2 x1431 0 u2 0 -1.34130711929499e-05
Rx1432 x1432 0 1
Fxc1432_1431 x1432 0 Vx1431 -158.15406128989
Cx1432 x1432 xm1432 1.01079656034734e-12
Vx1432 xm1432 0 0
Gx1432_2 x1432 0 u2 0 0.00212133168353545
Rx1433 x1433 0 1
Fxc1433_1434 x1433 0 Vx1434 3095.16001691797
Cx1433 x1433 xm1433 8.24832104280923e-14
Vx1433 xm1433 0 0
Gx1433_2 x1433 0 u2 0 -4.98084347666565e-08
Rx1434 x1434 0 1
Fxc1434_1433 x1434 0 Vx1433 -253.018034468733
Cx1434 x1434 xm1434 8.24832104280923e-14
Vx1434 xm1434 0 0
Gx1434_2 x1434 0 u2 0 1.26024322646235e-05
Rx1435 x1435 0 1
Fxc1435_1436 x1435 0 Vx1436 589.430233974696
Cx1435 x1435 xm1435 2.39433153810415e-13
Vx1435 xm1435 0 0
Gx1435_2 x1435 0 u2 0 -4.05529256563485e-07
Rx1436 x1436 0 1
Fxc1436_1435 x1436 0 Vx1435 -162.843855573984
Cx1436 x1436 xm1436 2.39433153810415e-13
Vx1436 xm1436 0 0
Gx1436_2 x1436 0 u2 0 6.60379476868495e-05
Rx1437 x1437 0 1
Fxc1437_1438 x1437 0 Vx1438 32.3873898502525
Cx1437 x1437 xm1437 2.46268600071512e-12
Vx1437 xm1437 0 0
Gx1437_2 x1437 0 u2 0 -0.00179486967652223
Rx1438 x1438 0 1
Fxc1438_1437 x1438 0 Vx1437 -31.8494183411198
Cx1438 x1438 xm1438 2.46268600071512e-12
Vx1438 xm1438 0 0
Gx1438_2 x1438 0 u2 0 0.0571655551953468
Rx1439 x1439 0 1
Fxc1439_1440 x1439 0 Vx1440 9.16604704249273
Cx1439 x1439 xm1439 3.96234308451514e-12
Vx1439 xm1439 0 0
Gx1439_2 x1439 0 u2 0 -0.000431172145165496
Rx1440 x1440 0 1
Fxc1440_1439 x1440 0 Vx1439 -55.494347398018
Cx1440 x1440 xm1440 3.96234308451514e-12
Vx1440 xm1440 0 0
Gx1440_2 x1440 0 u2 0 0.0239276168121626
Rx1441 x1441 0 1
Fxc1441_1442 x1441 0 Vx1442 208.578841102333
Cx1441 x1441 xm1441 8.60345839298812e-13
Vx1441 xm1441 0 0
Gx1441_2 x1441 0 u2 0 -3.62526071928876e-05
Rx1442 x1442 0 1
Fxc1442_1441 x1442 0 Vx1441 -38.2316422837127
Cx1442 x1442 xm1442 8.60345839298812e-13
Vx1442 xm1442 0 0
Gx1442_2 x1442 0 u2 0 0.00138599671005043
Rx1443 x1443 0 1
Fxc1443_1444 x1443 0 Vx1444 1269.74344070378
Cx1443 x1443 xm1443 9.68686303759719e-14
Vx1443 xm1443 0 0
Gx1443_2 x1443 0 u2 0 -1.95989950111513e-07
Rx1444 x1444 0 1
Fxc1444_1443 x1444 0 Vx1443 -493.64009076383
Cx1444 x1444 xm1444 9.68686303759719e-14
Vx1444 xm1444 0 0
Gx1444_2 x1444 0 u2 0 9.67484967618457e-05
Rx1445 x1445 0 1
Fxc1445_1446 x1445 0 Vx1446 57.6562075700509
Cx1445 x1445 xm1445 1.48715507116435e-12
Vx1445 xm1445 0 0
Gx1445_2 x1445 0 u2 0 -0.000348753086282661
Rx1446 x1446 0 1
Fxc1446_1445 x1446 0 Vx1445 -49.3815907808778
Cx1446 x1446 xm1446 1.48715507116435e-12
Vx1446 xm1446 0 0
Gx1446_2 x1446 0 u2 0 0.0172219821903785
Rx1447 x1447 0 1
Fxc1447_1448 x1447 0 Vx1448 122.987956973276
Cx1447 x1447 xm1447 4.21127124032637e-13
Vx1447 xm1447 0 0
Gx1447_2 x1447 0 u2 0 -1.30590329387355e-06
Rx1448 x1448 0 1
Fxc1448_1447 x1448 0 Vx1447 -294.477387037588
Cx1448 x1448 xm1448 4.21127124032637e-13
Vx1448 xm1448 0 0
Gx1448_2 x1448 0 u2 0 0.000384558989703662
Rx1449 x1449 0 1
Fxc1449_1450 x1449 0 Vx1450 770.371064458155
Cx1449 x1449 xm1449 2.74413394468355e-13
Vx1449 xm1449 0 0
Gx1449_2 x1449 0 u2 0 -4.22358911381612e-07
Rx1450 x1450 0 1
Fxc1450_1449 x1450 0 Vx1449 -117.319480514555
Cx1450 x1450 xm1450 2.74413394468355e-13
Vx1450 xm1450 0 0
Gx1450_2 x1450 0 u2 0 4.95509280739835e-05
Rx1451 x1451 0 1
Fxc1451_1452 x1451 0 Vx1452 37.0426242182526
Cx1451 x1451 xm1451 1.53173944244712e-12
Vx1451 xm1451 0 0
Gx1451_2 x1451 0 u2 0 -4.33040343427225e-05
Rx1452 x1452 0 1
Fxc1452_1451 x1452 0 Vx1451 -83.1008382816972
Cx1452 x1452 xm1452 1.53173944244712e-12
Vx1452 xm1452 0 0
Gx1452_2 x1452 0 u2 0 0.00359860155485964
Rx1453 x1453 0 1
Fxc1453_1454 x1453 0 Vx1454 5.72460876095774
Cx1453 x1453 xm1453 1.91528411913751e-13
Vx1453 xm1453 0 0
Gx1453_2 x1453 0 u2 0 -2.70165737945988e-09
Rx1454 x1454 0 1
Fxc1454_1453 x1454 0 Vx1453 -33446.4263272855
Cx1454 x1454 xm1454 1.91528411913751e-13
Vx1454 xm1454 0 0
Gx1454_2 x1454 0 u2 0 9.03607845036719e-05
Rx1455 x1455 0 1
Fxc1455_1456 x1455 0 Vx1456 1259.091033226
Cx1455 x1455 xm1455 2.36846187047956e-13
Vx1455 xm1455 0 0
Gx1455_2 x1455 0 u2 0 -2.71833957330908e-07
Rx1456 x1456 0 1
Fxc1456_1455 x1456 0 Vx1455 -119.830912068662
Cx1456 x1456 xm1456 2.36846187047956e-13
Vx1456 xm1456 0 0
Gx1456_2 x1456 0 u2 0 3.25741110381963e-05
Rx1457 x1457 0 1
Fxc1457_1458 x1457 0 Vx1458 36.0852726528186
Cx1457 x1457 xm1457 8.29948243480383e-13
Vx1457 xm1457 0 0
Gx1457_2 x1457 0 u2 0 -2.68051432615762e-06
Rx1458 x1458 0 1
Fxc1458_1457 x1458 0 Vx1457 -308.878497243482
Cx1458 x1458 xm1458 8.29948243480384e-13
Vx1458 xm1458 0 0
Gx1458_2 x1458 0 u2 0 0.000827953236903192
Rx1459 x1459 0 1
Fxc1459_1460 x1459 0 Vx1460 2124.5542048564
Cx1459 x1459 xm1459 1.49608073882079e-13
Vx1459 xm1459 0 0
Gx1459_2 x1459 0 u2 0 -1.54821120151765e-07
Rx1460 x1460 0 1
Fxc1460_1459 x1460 0 Vx1459 -154.566761679952
Cx1460 x1460 xm1460 1.49608073882079e-13
Vx1460 xm1460 0 0
Gx1460_2 x1460 0 u2 0 2.3930199181521e-05
Rx1461 x1461 0 1
Fxc1461_1462 x1461 0 Vx1462 232.279012952934
Cx1461 x1461 xm1461 8.78155428912643e-14
Vx1461 xm1461 0 0
Gx1461_2 x1461 0 u2 0 -1.16126006099731e-09
Rx1462 x1462 0 1
Fxc1462_1461 x1462 0 Vx1461 -4390.94147387229
Cx1462 x1462 xm1462 8.78155428912643e-14
Vx1462 xm1462 0 0
Gx1462_2 x1462 0 u2 0 5.09902496378456e-06
Rx1463 x1463 0 1
Fxc1463_1464 x1463 0 Vx1464 1478.76090862183
Cx1463 x1463 xm1463 4.67897291113138e-13
Vx1463 xm1463 0 0
Gx1463_2 x1463 0 u2 0 -4.89299708564559e-06
Rx1464 x1464 0 1
Fxc1464_1463 x1464 0 Vx1463 -19.0756792549105
Cx1464 x1464 xm1464 4.67897291113138e-13
Vx1464 xm1464 0 0
Gx1464_2 x1464 0 u2 0 9.33372430009871e-05
Rx1465 x1465 0 1
Fxc1465_1466 x1465 0 Vx1466 575.854584076211
Cx1465 x1465 xm1465 1.29257481425064e-13
Vx1465 xm1465 0 0
Gx1465_2 x1465 0 u2 0 -5.08176452576383e-08
Rx1466 x1466 0 1
Fxc1466_1465 x1466 0 Vx1465 -852.405821058812
Cx1466 x1466 xm1466 1.29257481425064e-13
Vx1466 xm1466 0 0
Gx1466_2 x1466 0 u2 0 4.33172566301127e-05
Rx1467 x1467 0 1
Fxc1467_1468 x1467 0 Vx1468 674.245588214102
Cx1467 x1467 xm1467 1.14664608873347e-13
Vx1467 xm1467 0 0
Gx1467_2 x1467 0 u2 0 -1.58551803856389e-07
Rx1468 x1468 0 1
Fxc1468_1467 x1468 0 Vx1467 -656.004705709629
Cx1468 x1468 xm1468 1.14664608873347e-13
Vx1468 xm1468 0 0
Gx1468_2 x1468 0 u2 0 0.000104010729428542
Rx1469 x1469 0 1
Fxc1469_1470 x1469 0 Vx1470 116.352316812739
Cx1469 x1469 xm1469 1.69186391030051e-12
Vx1469 xm1469 0 0
Gx1469_2 x1469 0 u2 0 -5.07139760509794e-05
Rx1470 x1470 0 1
Fxc1470_1469 x1470 0 Vx1469 -27.659160961593
Cx1470 x1470 xm1470 1.69186391030051e-12
Vx1470 xm1470 0 0
Gx1470_2 x1470 0 u2 0 0.00140270602659641
Rx1471 x1471 0 1
Fxc1471_1472 x1471 0 Vx1472 46.1458584356364
Cx1471 x1471 xm1471 5.92302008947924e-13
Vx1471 xm1471 0 0
Gx1471_2 x1471 0 u2 0 -7.00619715748342e-07
Rx1472 x1472 0 1
Fxc1472_1471 x1472 0 Vx1471 -582.112523305229
Cx1472 x1472 xm1472 5.92302008947924e-13
Vx1472 xm1472 0 0
Gx1472_2 x1472 0 u2 0 0.00040783951061166
Rx1473 x1473 0 1
Fxc1473_1474 x1473 0 Vx1474 13.4899120671812
Cx1473 x1473 xm1473 1.69585389952454e-11
Vx1473 xm1473 0 0
Gx1473_2 x1473 0 u2 0 -0.0657777436911043
Rx1474 x1474 0 1
Fxc1474_1473 x1474 0 Vx1473 -3.19889155237604
Cx1474 x1474 xm1474 1.69585389952454e-11
Vx1474 xm1474 0 0
Gx1474_2 x1474 0 u2 0 0.21041586862783
Rx1475 x1475 0 1
Fxc1475_1476 x1475 0 Vx1476 45.6455661572705
Cx1475 x1475 xm1475 2.98300305540713e-12
Vx1475 xm1475 0 0
Gx1475_2 x1475 0 u2 0 -0.000345280474005733
Rx1476 x1476 0 1
Fxc1476_1475 x1476 0 Vx1475 -28.1435898649539
Cx1476 x1476 xm1476 2.98300305540713e-12
Vx1476 xm1476 0 0
Gx1476_2 x1476 0 u2 0 0.00971743204879424
Rx1477 x1477 0 1
Fxc1477_1478 x1477 0 Vx1478 473.324234183567
Cx1477 x1477 xm1477 1.26171155346877e-12
Vx1477 xm1477 0 0
Gx1477_2 x1477 0 u2 0 -1.59187708051732e-05
Rx1478 x1478 0 1
Fxc1478_1477 x1478 0 Vx1477 -13.2361118145616
Cx1478 x1478 xm1478 1.26171155346877e-12
Vx1478 xm1478 0 0
Gx1478_2 x1478 0 u2 0 0.00021070263032765
Rx1479 x1479 0 1
Fxc1479_1480 x1479 0 Vx1480 35490.4690786351
Cx1479 x1479 xm1479 2.40296590857126e-13
Vx1479 xm1479 0 0
Gx1479_2 x1479 0 u2 0 -3.00930224402647e-07
Rx1480 x1480 0 1
Fxc1480_1479 x1480 0 Vx1479 -5.20509292560989
Cx1480 x1480 xm1480 2.40296590857126e-13
Vx1480 xm1480 0 0
Gx1480_2 x1480 0 u2 0 1.56636978214041e-06
Rx1481 x1481 0 1
Fxc1481_1482 x1481 0 Vx1482 375.437043371203
Cx1481 x1481 xm1481 7.07481712812474e-13
Vx1481 xm1481 0 0
Gx1481_2 x1481 0 u2 0 -3.43265494293932e-06
Rx1482 x1482 0 1
Fxc1482_1481 x1482 0 Vx1481 -58.0557529837625
Cx1482 x1482 xm1482 7.07481712812475e-13
Vx1482 xm1482 0 0
Gx1482_2 x1482 0 u2 0 0.000199285367445776
Rx1483 x1483 0 1
Fxc1483_1484 x1483 0 Vx1484 1.33655816675372
Cx1483 x1483 xm1483 2.47070341991198e-13
Vx1483 xm1483 0 0
Gx1483_2 x1483 0 u2 0 -4.65487670505573e-10
Rx1484 x1484 0 1
Fxc1484_1483 x1484 0 Vx1483 -123660.777440417
Cx1484 x1484 xm1484 2.47070341991198e-13
Vx1484 xm1484 0 0
Gx1484_2 x1484 0 u2 0 5.75625672236476e-05
Rx1485 x1485 0 1
Fxc1485_1486 x1485 0 Vx1486 643.678216101824
Cx1485 x1485 xm1485 6.42131520033378e-14
Vx1485 xm1485 0 0
Gx1485_2 x1485 0 u2 0 -7.97982611154097e-09
Rx1486 x1486 0 1
Fxc1486_1485 x1486 0 Vx1485 -3416.49935069765
Cx1486 x1486 xm1486 6.42131520033378e-14
Vx1486 xm1486 0 0
Gx1486_2 x1486 0 u2 0 2.72630707287599e-05
Rx1487 x1487 0 1
Fxc1487_1488 x1487 0 Vx1488 119.189992642376
Cx1487 x1487 xm1487 1.12198183373626e-11
Vx1487 xm1487 0 0
Gx1487_2 x1487 0 u2 0 -0.00196903726646598
Rx1488 x1488 0 1
Fxc1488_1487 x1488 0 Vx1487 -1.43502605193431
Cx1488 x1488 xm1488 1.12198183373626e-11
Vx1488 xm1488 0 0
Gx1488_2 x1488 0 u2 0 0.0028256197746082
Rx1489 x1489 0 1
Fxc1489_1490 x1489 0 Vx1490 3.74858034129987
Cx1489 x1489 xm1489 3.2472763080511e-12
Vx1489 xm1489 0 0
Gx1489_2 x1489 0 u2 0 -6.86976422616017e-05
Rx1490 x1490 0 1
Fxc1490_1489 x1490 0 Vx1489 -307.099474521271
Cx1490 x1490 xm1490 3.2472763080511e-12
Vx1490 xm1490 0 0
Gx1490_2 x1490 0 u2 0 0.0210970098393882
Rx1491 x1491 0 1
Fxc1491_1492 x1491 0 Vx1492 5.28329475425347
Cx1491 x1491 xm1491 3.71285809172693e-12
Vx1491 xm1491 0 0
Gx1491_2 x1491 0 u2 0 -6.55879280884544e-05
Rx1492 x1492 0 1
Fxc1492_1491 x1492 0 Vx1491 -182.502201406073
Cx1492 x1492 xm1492 3.71285809172693e-12
Vx1492 xm1492 0 0
Gx1492_2 x1492 0 u2 0 0.0119699412618061
Rx1493 x1493 0 1
Fxc1493_1494 x1493 0 Vx1494 6.3409246812571
Cx1493 x1493 xm1493 7.59177081056463e-13
Vx1493 xm1493 0 0
Gx1493_2 x1493 0 u2 0 -1.43389071404067e-07
Rx1494 x1494 0 1
Fxc1494_1493 x1494 0 Vx1493 -3492.5454298433
Cx1494 x1494 xm1494 7.59177081056463e-13
Vx1494 xm1494 0 0
Gx1494_2 x1494 0 u2 0 0.00050079284602175
Rx1495 x1495 0 1
Fxc1495_1496 x1495 0 Vx1496 230.643356966458
Cx1495 x1495 xm1495 2.02585528546519e-13
Vx1495 xm1495 0 0
Gx1495_2 x1495 0 u2 0 -1.04286172096209e-07
Rx1496 x1496 0 1
Fxc1496_1495 x1496 0 Vx1495 -1292.73472729722
Cx1496 x1496 xm1496 2.02585528546519e-13
Vx1496 xm1496 0 0
Gx1496_2 x1496 0 u2 0 0.000134814356245663
Rx1497 x1497 0 1
Fxc1497_1498 x1497 0 Vx1498 724.974623088263
Cx1497 x1497 xm1497 4.24372223574733e-14
Vx1497 xm1497 0 0
Gx1497_2 x1497 0 u2 0 -7.06216793609314e-09
Rx1498 x1498 0 1
Fxc1498_1497 x1498 0 Vx1497 -10407.4965125006
Cx1498 x1498 xm1498 4.24372223574733e-14
Vx1498 xm1498 0 0
Gx1498_2 x1498 0 u2 0 7.34994881655831e-05
Rx1499 x1499 0 1
Fxc1499_1500 x1499 0 Vx1500 1475.40988353595
Cx1499 x1499 xm1499 1.00885100580125e-13
Vx1499 xm1499 0 0
Gx1499_2 x1499 0 u2 0 -6.04980876332292e-08
Rx1500 x1500 0 1
Fxc1500_1499 x1500 0 Vx1499 -972.781125520802
Cx1500 x1500 xm1500 1.00885100580125e-13
Vx1500 xm1500 0 0
Gx1500_2 x1500 0 u2 0 5.88513977797089e-05
Rx1501 x1501 0 1
Fxc1501_1502 x1501 0 Vx1502 125.413451486806
Cx1501 x1501 xm1501 4.00195036079336e-13
Vx1501 xm1501 0 0
Gx1501_2 x1501 0 u2 0 -3.31391916706323e-07
Rx1502 x1502 0 1
Fxc1502_1501 x1502 0 Vx1501 -580.792504414272
Cx1502 x1502 xm1502 4.00195036079336e-13
Vx1502 xm1502 0 0
Gx1502_2 x1502 0 u2 0 0.000192469941246511
Rx1503 x1503 0 1
Fxc1503_1504 x1503 0 Vx1504 9.56568027582822
Cx1503 x1503 xm1503 2.78329702880848e-13
Vx1503 xm1503 0 0
Gx1503_2 x1503 0 u2 0 -5.53563934265562e-09
Rx1504 x1504 0 1
Fxc1504_1503 x1504 0 Vx1503 -20508.6895623213
Cx1504 x1504 xm1504 2.78329702880848e-13
Vx1504 xm1504 0 0
Gx1504_2 x1504 0 u2 0 0.000113528708807497
Rx1505 x1505 0 1
Fxc1505_1506 x1505 0 Vx1506 62.3715380064075
Cx1505 x1505 xm1505 1.59370707888504e-12
Vx1505 xm1505 0 0
Gx1505_2 x1505 0 u2 0 -1.43857389269971e-05
Rx1506 x1506 0 1
Fxc1506_1505 x1506 0 Vx1505 -106.192728825299
Cx1506 x1506 xm1506 1.59370707888504e-12
Vx1506 xm1506 0 0
Gx1506_2 x1506 0 u2 0 0.00152766087282615
Rx1507 x1507 0 1
Fxc1507_1508 x1507 0 Vx1508 229.689184071515
Cx1507 x1507 xm1507 1.50328460311422e-12
Vx1507 xm1507 0 0
Gx1507_2 x1507 0 u2 0 -1.65311083485886e-05
Rx1508 x1508 0 1
Fxc1508_1507 x1508 0 Vx1507 -34.1916165399867
Cx1508 x1508 xm1508 1.50328460311422e-12
Vx1508 xm1508 0 0
Gx1508_2 x1508 0 u2 0 0.000565225317635916
Rx1509 x1509 0 1
Fxc1509_1510 x1509 0 Vx1510 96.6589763152531
Cx1509 x1509 xm1509 2.99713440633919e-12
Vx1509 xm1509 0 0
Gx1509_2 x1509 0 u2 0 -0.000147932228049142
Rx1510 x1510 0 1
Fxc1510_1509 x1510 0 Vx1509 -19.0085566528686
Cx1510 x1510 xm1510 2.99713440633919e-12
Vx1510 xm1510 0 0
Gx1510_2 x1510 0 u2 0 0.0028119781376572
Rx1511 x1511 0 1
Fxc1511_1512 x1511 0 Vx1512 13201.8644241837
Cx1511 x1511 xm1511 4.59729955117924e-13
Vx1511 xm1511 0 0
Gx1511_2 x1511 0 u2 0 -3.39969344570208e-07
Rx1512 x1512 0 1
Fxc1512_1511 x1512 0 Vx1511 -5.65310352397753
Cx1512 x1512 xm1512 4.59729955117924e-13
Vx1512 xm1512 0 0
Gx1512_2 x1512 0 u2 0 1.92188189983417e-06
Rx1513 x1513 0 1
Fxc1513_1514 x1513 0 Vx1514 5.67131389681892
Cx1513 x1513 xm1513 2.42031501813512e-12
Vx1513 xm1513 0 0
Gx1513_2 x1513 0 u2 0 -6.38305096899387e-06
Rx1514 x1514 0 1
Fxc1514_1513 x1514 0 Vx1513 -547.020496816947
Cx1514 x1514 xm1514 2.42031501813512e-12
Vx1514 xm1514 0 0
Gx1514_2 x1514 0 u2 0 0.00349165971226692
Rx1515 x1515 0 1
Fxc1515_1516 x1515 0 Vx1516 63.2648897001453
Cx1515 x1515 xm1515 5.54877528405509e-13
Vx1515 xm1515 0 0
Gx1515_2 x1515 0 u2 0 -1.53421681408806e-07
Rx1516 x1516 0 1
Fxc1516_1515 x1516 0 Vx1515 -984.345304088486
Cx1516 x1516 xm1516 5.54877528405509e-13
Vx1516 xm1516 0 0
Gx1516_2 x1516 0 u2 0 0.000151019911640118
Rx1517 x1517 0 1
Cx1517 x1517 0 1.61089900076846e-09
Gx1517_2 x1517 0 u2 0 -1.59809499057346
Rx1518 x1518 0 1
Fxc1518_1519 x1518 0 Vx1519 1.10283582237019
Cx1518 x1518 xm1518 2.19812424587013e-10
Vx1518 xm1518 0 0
Gx1518_2 x1518 0 u2 0 -0.0733580247132006
Rx1519 x1519 0 1
Fxc1519_1518 x1519 0 Vx1518 -7.67587001499757
Cx1519 x1519 xm1519 2.19812424587013e-10
Vx1519 xm1519 0 0
Gx1519_2 x1519 0 u2 0 0.563086662255507
Rx1520 x1520 0 1
Fxc1520_1521 x1520 0 Vx1521 6.35136205952906
Cx1520 x1520 xm1520 1.87705184078918e-09
Vx1520 xm1520 0 0
Gx1520_2 x1520 0 u2 0 -0.313428114236027
Rx1521 x1521 0 1
Fxc1521_1520 x1521 0 Vx1520 -0.191940354015187
Cx1521 x1521 xm1521 1.87705184078918e-09
Vx1521 xm1521 0 0
Gx1521_2 x1521 0 u2 0 0.0601595032047757
Rx1522 x1522 0 1
Fxc1522_1523 x1522 0 Vx1523 3.95959125789346
Cx1522 x1522 xm1522 4.32510417049148e-11
Vx1522 xm1522 0 0
Gx1522_2 x1522 0 u2 0 -3.96060512552686e-06
Rx1523 x1523 0 1
Fxc1523_1522 x1523 0 Vx1522 -304.117346171678
Cx1523 x1523 xm1523 4.32510417049148e-11
Vx1523 xm1523 0 0
Gx1523_2 x1523 0 u2 0 0.00120448872000918
Rx1524 x1524 0 1
Fxc1524_1525 x1524 0 Vx1525 196.048665379505
Cx1524 x1524 xm1524 6.12250410889856e-12
Vx1524 xm1524 0 0
Gx1524_2 x1524 0 u2 0 -3.38878735837355e-06
Rx1525 x1525 0 1
Fxc1525_1524 x1525 0 Vx1524 -150.276850665396
Cx1525 x1525 xm1525 6.12250410889856e-12
Vx1525 xm1525 0 0
Gx1525_2 x1525 0 u2 0 0.000509256291791084
Rx1526 x1526 0 1
Fxc1526_1527 x1526 0 Vx1527 126.258049380707
Cx1526 x1526 xm1526 4.14799482577559e-11
Vx1526 xm1526 0 0
Gx1526_2 x1526 0 u2 0 -0.0273566650336182
Rx1527 x1527 0 1
Fxc1527_1526 x1527 0 Vx1526 -0.250997317312743
Cx1527 x1527 xm1527 4.14799482577559e-11
Vx1527 xm1527 0 0
Gx1527_2 x1527 0 u2 0 0.0068664495340615
Rx1528 x1528 0 1
Fxc1528_1529 x1528 0 Vx1529 21988.3340192612
Cx1528 x1528 xm1528 1.45549226115441e-14
Vx1528 xm1528 0 0
Gx1528_2 x1528 0 u2 0 -3.27122049462339e-09
Rx1529 x1529 0 1
Fxc1529_1528 x1529 0 Vx1528 -4411.50704730986
Cx1529 x1529 xm1529 1.45549226115441e-14
Vx1529 xm1529 0 0
Gx1529_2 x1529 0 u2 0 1.44310122653355e-05
Rx1530 x1530 0 1
Fxc1530_1531 x1530 0 Vx1531 21.1331721863719
Cx1530 x1530 xm1530 1.60409482204103e-11
Vx1530 xm1530 0 0
Gx1530_2 x1530 0 u2 0 -0.00214748036831327
Rx1531 x1531 0 1
Fxc1531_1530 x1531 0 Vx1530 -6.56793525804424
Cx1531 x1531 xm1531 1.60409482204103e-11
Vx1531 xm1531 0 0
Gx1531_2 x1531 0 u2 0 0.0141045120270026
Rx1532 x1532 0 1
Fxc1532_1533 x1532 0 Vx1533 5.95881996256681
Cx1532 x1532 xm1532 1.87789127101595e-11
Vx1532 xm1532 0 0
Gx1532_2 x1532 0 u2 0 -0.000683844520376207
Rx1533 x1533 0 1
Fxc1533_1532 x1533 0 Vx1532 -36.4130839798716
Cx1533 x1533 xm1533 1.87789127101595e-11
Vx1533 xm1533 0 0
Gx1533_2 x1533 0 u2 0 0.0249008879496338
Rx1534 x1534 0 1
Fxc1534_1535 x1534 0 Vx1535 58.0726784354013
Cx1534 x1534 xm1534 1.4701859252872e-12
Vx1534 xm1534 0 0
Gx1534_2 x1534 0 u2 0 -1.71997301236869e-06
Rx1535 x1535 0 1
Fxc1535_1534 x1535 0 Vx1534 -209.574292792984
Cx1535 x1535 xm1535 1.4701859252872e-12
Vx1535 xm1535 0 0
Gx1535_2 x1535 0 u2 0 0.000360462127690187
Rx1536 x1536 0 1
Fxc1536_1537 x1536 0 Vx1537 256.305706779398
Cx1536 x1536 xm1536 2.39937551270491e-13
Vx1536 xm1536 0 0
Gx1536_2 x1536 0 u2 0 -2.13033982736333e-08
Rx1537 x1537 0 1
Fxc1537_1536 x1537 0 Vx1536 -1526.19260674663
Cx1537 x1537 xm1537 2.39937551270491e-13
Vx1537 xm1537 0 0
Gx1537_2 x1537 0 u2 0 3.2513088943798e-05
Rx1538 x1538 0 1
Fxc1538_1539 x1538 0 Vx1539 713.834655162133
Cx1538 x1538 xm1538 3.58178612159909e-13
Vx1538 xm1538 0 0
Gx1538_2 x1538 0 u2 0 -1.4540286333917e-07
Rx1539 x1539 0 1
Fxc1539_1538 x1539 0 Vx1538 -299.925406894304
Cx1539 x1539 xm1539 3.58178612159909e-13
Vx1539 xm1539 0 0
Gx1539_2 x1539 0 u2 0 4.36100129505975e-05
Rx1540 x1540 0 1
Fxc1540_1541 x1540 0 Vx1541 39.2639489169957
Cx1540 x1540 xm1540 5.21591991919758e-12
Vx1540 xm1540 0 0
Gx1540_2 x1540 0 u2 0 -6.49101452816451e-05
Rx1541 x1541 0 1
Fxc1541_1540 x1541 0 Vx1540 -67.2978726905257
Cx1541 x1541 xm1541 5.21591991919758e-12
Vx1541 xm1541 0 0
Gx1541_2 x1541 0 u2 0 0.00436831469348768
Rx1542 x1542 0 1
Fxc1542_1543 x1542 0 Vx1543 35.3646991426765
Cx1542 x1542 xm1542 9.36281020722465e-13
Vx1542 xm1542 0 0
Gx1542_2 x1542 0 u2 0 -3.22841542421718e-07
Rx1543 x1543 0 1
Fxc1543_1542 x1543 0 Vx1542 -763.619337219721
Cx1543 x1543 xm1543 9.36281020722465e-13
Vx1543 xm1543 0 0
Gx1543_2 x1543 0 u2 0 0.000246528044651064
Rx1544 x1544 0 1
Fxc1544_1545 x1544 0 Vx1545 221.526299864096
Cx1544 x1544 xm1544 5.00909331659054e-13
Vx1544 xm1544 0 0
Gx1544_2 x1544 0 u2 0 -5.12521701462589e-08
Rx1545 x1545 0 1
Fxc1545_1544 x1545 0 Vx1544 -1089.2087144039
Cx1545 x1545 xm1545 5.00909331659054e-13
Vx1545 xm1545 0 0
Gx1545_2 x1545 0 u2 0 5.58243103554167e-05
Rx1546 x1546 0 1
Fxc1546_1547 x1546 0 Vx1547 334.906543793632
Cx1546 x1546 xm1546 2.21603934379445e-12
Vx1546 xm1546 0 0
Gx1546_2 x1546 0 u2 0 -4.38909788905065e-06
Rx1547 x1547 0 1
Fxc1547_1546 x1547 0 Vx1546 -29.2237485470108
Cx1547 x1547 xm1547 2.21603934379444e-12
Vx1547 xm1547 0 0
Gx1547_2 x1547 0 u2 0 0.000128265893057832
Rx1548 x1548 0 1
Fxc1548_1549 x1548 0 Vx1549 17001.6380250491
Cx1548 x1548 xm1548 1.03257318571619e-14
Vx1548 xm1548 0 0
Gx1548_2 x1548 0 u2 0 -2.94122800405986e-09
Rx1549 x1549 0 1
Fxc1549_1548 x1549 0 Vx1548 -18232.7304267604
Cx1549 x1549 xm1549 1.03257318571619e-14
Vx1549 xm1549 0 0
Gx1549_2 x1549 0 u2 0 5.3626617321662e-05
Rx1550 x1550 0 1
Fxc1550_1551 x1550 0 Vx1551 7580.63241325557
Cx1550 x1550 xm1550 2.74819843338129e-12
Vx1550 xm1550 0 0
Gx1550_2 x1550 0 u2 0 -2.6202833316178e-05
Rx1551 x1551 0 1
Fxc1551_1550 x1551 0 Vx1550 -0.527297167993212
Cx1551 x1551 xm1551 2.74819843338129e-12
Vx1551 xm1551 0 0
Gx1551_2 x1551 0 u2 0 1.38166798010188e-05
Rx1552 x1552 0 1
Fxc1552_1553 x1552 0 Vx1553 330.150555703687
Cx1552 x1552 xm1552 4.24036342517206e-12
Vx1552 xm1552 0 0
Gx1552_2 x1552 0 u2 0 -2.7798048785484e-05
Rx1553 x1553 0 1
Fxc1553_1552 x1553 0 Vx1552 -7.52849052181352
Cx1553 x1553 xm1553 4.24036342517206e-12
Vx1553 xm1553 0 0
Gx1553_2 x1553 0 u2 0 0.000209277346806426
Rx1554 x1554 0 1
Fxc1554_1555 x1554 0 Vx1555 1164.26845642317
Cx1554 x1554 xm1554 9.58496587203372e-13
Vx1554 xm1554 0 0
Gx1554_2 x1554 0 u2 0 -9.85355298544214e-07
Rx1555 x1555 0 1
Fxc1555_1554 x1555 0 Vx1554 -38.8974643800463
Cx1555 x1555 xm1555 9.58496587203372e-13
Vx1555 xm1555 0 0
Gx1555_2 x1555 0 u2 0 3.83278226268134e-05
Rx1556 x1556 0 1
Fxc1556_1557 x1556 0 Vx1557 213.451660276106
Cx1556 x1556 xm1556 1.12815467078128e-12
Vx1556 xm1556 0 0
Gx1556_2 x1556 0 u2 0 -1.12307780104608e-06
Rx1557 x1557 0 1
Fxc1557_1556 x1557 0 Vx1556 -131.831523950433
Cx1557 x1557 xm1557 1.12815467078128e-12
Vx1557 xm1557 0 0
Gx1557_2 x1557 0 u2 0 0.000148057058026806
Rx1558 x1558 0 1
Fxc1558_1559 x1558 0 Vx1559 32.8263627611749
Cx1558 x1558 xm1558 1.79517864865178e-12
Vx1558 xm1558 0 0
Gx1558_2 x1558 0 u2 0 -2.70905999901583e-06
Rx1559 x1559 0 1
Fxc1559_1558 x1559 0 Vx1558 -291.318109924474
Cx1559 x1559 xm1559 1.79517864865178e-12
Vx1559 xm1559 0 0
Gx1559_2 x1559 0 u2 0 0.000789198238585289
Rx1560 x1560 0 1
Fxc1560_1561 x1560 0 Vx1561 679.734283805673
Cx1560 x1560 xm1560 6.11941306890275e-13
Vx1560 xm1560 0 0
Gx1560_2 x1560 0 u2 0 -4.33716700256784e-07
Rx1561 x1561 0 1
Fxc1561_1560 x1561 0 Vx1560 -91.2380382457165
Cx1561 x1561 xm1561 6.11941306890275e-13
Vx1561 xm1561 0 0
Gx1561_2 x1561 0 u2 0 3.95714608858345e-05
Rx1562 x1562 0 1
Fxc1562_1563 x1562 0 Vx1563 56.6817645759923
Cx1562 x1562 xm1562 1.42015889054634e-12
Vx1562 xm1562 0 0
Gx1562_2 x1562 0 u2 0 -5.33614901713773e-07
Rx1563 x1563 0 1
Fxc1563_1562 x1563 0 Vx1562 -466.817505667653
Cx1563 x1563 xm1563 1.42015889054634e-12
Vx1563 xm1563 0 0
Gx1563_2 x1563 0 u2 0 0.000249100777405113
Rx1564 x1564 0 1
Fxc1564_1565 x1564 0 Vx1565 34.9090735740061
Cx1564 x1564 xm1564 7.91863406834521e-12
Vx1564 xm1564 0 0
Gx1564_2 x1564 0 u2 0 -0.00029570848248748
Rx1565 x1565 0 1
Fxc1565_1564 x1565 0 Vx1564 -32.7802160498318
Cx1565 x1565 xm1565 7.91863406834521e-12
Vx1565 xm1565 0 0
Gx1565_2 x1565 0 u2 0 0.00969338794370752
Rx1566 x1566 0 1
Fxc1566_1567 x1566 0 Vx1567 849.912088117841
Cx1566 x1566 xm1566 9.12011682999143e-13
Vx1566 xm1566 0 0
Gx1566_2 x1566 0 u2 0 -3.59703092665933e-07
Rx1567 x1567 0 1
Fxc1567_1566 x1567 0 Vx1566 -119.585984142478
Cx1567 x1567 xm1567 9.12011682999143e-13
Vx1567 xm1567 0 0
Gx1567_2 x1567 0 u2 0 4.30154483355484e-05
Rx1568 x1568 0 1
Fxc1568_1569 x1568 0 Vx1569 101.147868350739
Cx1568 x1568 xm1568 2.64454642404486e-12
Vx1568 xm1568 0 0
Gx1568_2 x1568 0 u2 0 -1.65992107672464e-06
Rx1569 x1569 0 1
Fxc1569_1568 x1569 0 Vx1568 -132.271577310423
Cx1569 x1569 xm1569 2.64454642404486e-12
Vx1569 xm1569 0 0
Gx1569_2 x1569 0 u2 0 0.000219560379029185
Rx1570 x1570 0 1
Fxc1570_1571 x1570 0 Vx1571 33.2593824265232
Cx1570 x1570 xm1570 1.51286572624691e-11
Vx1570 xm1570 0 0
Gx1570_2 x1570 0 u2 0 -0.000186582528054369
Rx1571 x1571 0 1
Fxc1571_1570 x1571 0 Vx1570 -17.6646694676801
Cx1571 x1571 xm1571 1.51286572624691e-11
Vx1571 xm1571 0 0
Gx1571_2 x1571 0 u2 0 0.00329591868652459
Rx1572 x1572 0 1
Fxc1572_1573 x1572 0 Vx1573 3.87336369442715
Cx1572 x1572 xm1572 1.22419165937248e-10
Vx1572 xm1572 0 0
Gx1572_2 x1572 0 u2 0 -0.0362447013326694
Rx1573 x1573 0 1
Fxc1573_1572 x1573 0 Vx1572 -5.42872386522244
Cx1573 x1573 xm1573 1.22419165937248e-10
Vx1573 xm1573 0 0
Gx1573_2 x1573 0 u2 0 0.196762475112522
Rx1574 x1574 0 1
Fxc1574_1575 x1574 0 Vx1575 143.460527178785
Cx1574 x1574 xm1574 1.76967136661136e-11
Vx1574 xm1574 0 0
Gx1574_2 x1574 0 u2 0 -9.6455488452902e-05
Rx1575 x1575 0 1
Fxc1575_1574 x1575 0 Vx1574 -4.73046350824725
Cx1575 x1575 xm1575 1.76967136661136e-11
Vx1575 xm1575 0 0
Gx1575_2 x1575 0 u2 0 0.000456279168296618
Rx1576 x1576 0 1
Fxc1576_1577 x1576 0 Vx1577 2.01557203114741
Cx1576 x1576 xm1576 1.26800162802138e-11
Vx1576 xm1576 0 0
Gx1576_2 x1576 0 u2 0 -1.37559224793841e-06
Rx1577 x1577 0 1
Fxc1577_1576 x1577 0 Vx1576 -794.198370559574
Cx1577 x1577 xm1577 1.26800162802138e-11
Vx1577 xm1577 0 0
Gx1577_2 x1577 0 u2 0 0.00109249312186707
Rx1578 x1578 0 1
Cx1578 x1578 0 7.05227504597918e-09
Gx1578_2 x1578 0 u2 0 -1.69557023065726
Rx1579 x1579 0 1
Fxc1579_1580 x1579 0 Vx1580 225.728703794371
Cx1579 x1579 xm1579 1.15460286288366e-12
Vx1579 xm1579 0 0
Gx1579_2 x1579 0 u2 0 -9.58180319929274e-07
Rx1580 x1580 0 1
Fxc1580_1579 x1580 0 Vx1579 -127.578343173863
Cx1580 x1580 xm1580 1.15460286288366e-12
Vx1580 xm1580 0 0
Gx1580_2 x1580 0 u2 0 0.000122243057678379
Rx1581 x1581 0 1
Fxc1581_1582 x1581 0 Vx1582 9.05504448124067
Cx1581 x1581 xm1581 2.18132271178657e-10
Vx1581 xm1581 0 0
Gx1581_2 x1581 0 u2 0 -9.73091817660008e-05
Rx1582 x1582 0 1
Fxc1582_1581 x1582 0 Vx1581 -35.7098077712971
Cx1582 x1582 xm1582 2.18132271178657e-10
Vx1582 xm1582 0 0
Gx1582_2 x1582 0 u2 0 0.0034748921752461
Rx1583 x1583 0 1
Fxc1583_1584 x1583 0 Vx1584 7.42699481325217
Cx1583 x1583 xm1583 8.40037698819289e-11
Vx1583 xm1583 0 0
Gx1583_2 x1583 0 u2 0 -0.00449698915680542
Rx1584 x1584 0 1
Fxc1584_1583 x1584 0 Vx1583 -8.91756035539826
Cx1584 x1584 xm1584 8.40037698819289e-11
Vx1584 xm1584 0 0
Gx1584_2 x1584 0 u2 0 0.0401021722233839
Rx1585 x1585 0 1
Fxc1585_1586 x1585 0 Vx1586 6.76257349855225
Cx1585 x1585 xm1585 5.30998399535694e-11
Vx1585 xm1585 0 0
Gx1585_2 x1585 0 u2 0 -0.000117804816363985
Rx1586 x1586 0 1
Fxc1586_1585 x1586 0 Vx1585 -36.2370460750124
Cx1586 x1586 xm1586 5.30998399535694e-11
Vx1586 xm1586 0 0
Gx1586_2 x1586 0 u2 0 0.00426889855844009
Rx1587 x1587 0 1
Fxc1587_1588 x1587 0 Vx1588 239.140501229814
Cx1587 x1587 xm1587 1.35912169198298e-12
Vx1587 xm1587 0 0
Gx1587_2 x1587 0 u2 0 -3.62388784840492e-07
Rx1588 x1588 0 1
Fxc1588_1587 x1588 0 Vx1587 -229.745159069808
Cx1588 x1588 xm1588 1.35912169198298e-12
Vx1588 xm1588 0 0
Gx1588_2 x1588 0 u2 0 8.32570690182933e-05
Rx1589 x1589 0 1
Fxc1589_1590 x1589 0 Vx1590 43.2013103157405
Cx1589 x1589 xm1589 6.31264225400471e-12
Vx1589 xm1589 0 0
Gx1589_2 x1589 0 u2 0 -1.1637928145185e-05
Rx1590 x1590 0 1
Fxc1590_1589 x1590 0 Vx1589 -63.8606713142529
Cx1590 x1590 xm1590 6.31264225400471e-12
Vx1590 xm1590 0 0
Gx1590_2 x1590 0 u2 0 0.000743205904058555
Rx1591 x1591 0 1
Fxc1591_1592 x1591 0 Vx1592 0.867802741268697
Cx1591 x1591 xm1591 1.33436643953763e-11
Vx1591 xm1591 0 0
Gx1591_2 x1591 0 u2 0 -7.48318242340968e-06
Rx1592 x1592 0 1
Fxc1592_1591 x1592 0 Vx1591 -963.364418640562
Cx1592 x1592 xm1592 1.33436643953763e-11
Vx1592 xm1592 0 0
Gx1592_2 x1592 0 u2 0 0.00720903168490934
Rx1593 x1593 0 1
Fxc1593_1594 x1593 0 Vx1594 216.701203294362
Cx1593 x1593 xm1593 1.32642627349223e-11
Vx1593 xm1593 0 0
Gx1593_2 x1593 0 u2 0 -2.38956196572277e-05
Rx1594 x1594 0 1
Fxc1594_1593 x1594 0 Vx1593 -8.07337773373533
Cx1594 x1594 xm1594 1.32642627349223e-11
Vx1594 xm1594 0 0
Gx1594_2 x1594 0 u2 0 0.00019291836367447
Rx1595 x1595 0 1
Fxc1595_1596 x1595 0 Vx1596 19.7129407412976
Cx1595 x1595 xm1595 1.08698420955425e-11
Vx1595 xm1595 0 0
Gx1595_2 x1595 0 u2 0 -1.76812595167102e-05
Rx1596 x1596 0 1
Fxc1596_1595 x1596 0 Vx1595 -76.1607475176606
Cx1596 x1596 xm1596 1.08698420955425e-11
Vx1596 xm1596 0 0
Gx1596_2 x1596 0 u2 0 0.0013466179418464
Rx1597 x1597 0 1
Fxc1597_1598 x1597 0 Vx1598 92.685475334831
Cx1597 x1597 xm1597 4.56998680318091e-12
Vx1597 xm1597 0 0
Gx1597_2 x1597 0 u2 0 -9.45003185010707e-06
Rx1598 x1598 0 1
Fxc1598_1597 x1598 0 Vx1597 -78.9965325420085
Cx1598 x1598 xm1598 4.56998680318091e-12
Vx1598 xm1598 0 0
Gx1598_2 x1598 0 u2 0 0.00074651974857
Rx1599 x1599 0 1
Cx1599 x1599 0 1.02081938428761e-08
Gx1599_2 x1599 0 u2 0 -1.29426055272561
Rx1600 x1600 0 1
Fxc1600_1601 x1600 0 Vx1601 18.8021931553848
Cx1600 x1600 xm1600 1.53254609092949e-11
Vx1600 xm1600 0 0
Gx1600_2 x1600 0 u2 0 -1.46157699240128e-05
Rx1601 x1601 0 1
Fxc1601_1600 x1601 0 Vx1600 -96.9359611002553
Cx1601 x1601 xm1601 1.53254609092949e-11
Vx1601 xm1601 0 0
Gx1601_2 x1601 0 u2 0 0.00141679370480439
Rx1602 x1602 0 1
Cx1602 x1602 0 5.04506053260489e-08
Gx1602_2 x1602 0 u2 0 -0.55208238084925
Gyc1_1 y1 0 x1 0 -1
Gyc1_2 y1 0 x2 0 1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 -1
Gyc1_6 y1 0 x6 0 1
Gyc1_7 y1 0 x7 0 1
Gyc1_8 y1 0 x8 0 -1
Gyc1_9 y1 0 x9 0 1
Gyc1_10 y1 0 x10 0 -1
Gyc1_11 y1 0 x11 0 1
Gyc1_12 y1 0 x12 0 -1
Gyc1_13 y1 0 x13 0 -1
Gyc1_14 y1 0 x14 0 1
Gyc1_15 y1 0 x15 0 1
Gyc1_16 y1 0 x16 0 1
Gyc1_17 y1 0 x17 0 -1
Gyc1_18 y1 0 x18 0 1
Gyc1_19 y1 0 x19 0 1
Gyc1_20 y1 0 x20 0 1
Gyc1_21 y1 0 x21 0 -1
Gyc1_22 y1 0 x22 0 -1
Gyc1_23 y1 0 x23 0 -1
Gyc1_24 y1 0 x24 0 1
Gyc1_25 y1 0 x25 0 -1
Gyc1_26 y1 0 x26 0 1
Gyc1_27 y1 0 x27 0 -1
Gyc1_28 y1 0 x28 0 1
Gyc1_29 y1 0 x29 0 -1
Gyc1_30 y1 0 x30 0 1
Gyc1_31 y1 0 x31 0 -1
Gyc1_32 y1 0 x32 0 1
Gyc1_33 y1 0 x33 0 -1
Gyc1_34 y1 0 x34 0 1
Gyc1_35 y1 0 x35 0 -1
Gyc1_36 y1 0 x36 0 -1
Gyc1_37 y1 0 x37 0 1
Gyc1_38 y1 0 x38 0 -1
Gyc1_39 y1 0 x39 0 1
Gyc1_40 y1 0 x40 0 0.562823070074008
Gyc1_41 y1 0 x41 0 -1
Gyc1_42 y1 0 x42 0 1
Gyc1_43 y1 0 x43 0 1
Gyc1_44 y1 0 x44 0 1
Gyc1_45 y1 0 x45 0 -1
Gyc1_46 y1 0 x46 0 1
Gyc1_47 y1 0 x47 0 -1
Gyc1_48 y1 0 x48 0 -1
Gyc1_49 y1 0 x49 0 1
Gyc1_50 y1 0 x50 0 1
Gyc1_51 y1 0 x51 0 1
Gyc1_52 y1 0 x52 0 1
Gyc1_53 y1 0 x53 0 -1
Gyc1_54 y1 0 x54 0 1
Gyc1_55 y1 0 x55 0 -1
Gyc1_56 y1 0 x56 0 1
Gyc1_57 y1 0 x57 0 1
Gyc1_58 y1 0 x58 0 -1
Gyc1_59 y1 0 x59 0 -1
Gyc1_60 y1 0 x60 0 -1
Gyc1_61 y1 0 x61 0 0.706400192735412
Gyc1_62 y1 0 x62 0 -1
Gyc1_63 y1 0 x63 0 1
Gyc1_64 y1 0 x64 0 1
Gyc1_65 y1 0 x65 0 1
Gyc1_66 y1 0 x66 0 1
Gyc1_67 y1 0 x67 0 -1
Gyc1_68 y1 0 x68 0 1
Gyc1_69 y1 0 x69 0 -1
Gyc1_70 y1 0 x70 0 -1
Gyc1_71 y1 0 x71 0 -1
Gyc1_72 y1 0 x72 0 -1
Gyc1_73 y1 0 x73 0 1
Gyc1_74 y1 0 x74 0 -1
Gyc1_75 y1 0 x75 0 -1
Gyc1_76 y1 0 x76 0 -1
Gyc1_77 y1 0 x77 0 1
Gyc1_78 y1 0 x78 0 1
Gyc1_79 y1 0 x79 0 -1
Gyc1_80 y1 0 x80 0 1
Gyc1_81 y1 0 x81 0 1
Gyc1_82 y1 0 x82 0 -1
Gyc1_83 y1 0 x83 0 -1
Gyc1_84 y1 0 x84 0 -1
Gyc1_85 y1 0 x85 0 1
Gyc1_86 y1 0 x86 0 1
Gyc1_87 y1 0 x87 0 -1
Gyc1_88 y1 0 x88 0 -1
Gyc1_89 y1 0 x89 0 1
Gyc1_90 y1 0 x90 0 -1
Gyc1_91 y1 0 x91 0 1
Gyc1_92 y1 0 x92 0 -0.190381393765198
Gyc1_93 y1 0 x93 0 1
Gyc1_94 y1 0 x94 0 -1
Gyc1_95 y1 0 x95 0 -1
Gyc1_96 y1 0 x96 0 -1
Gyc1_97 y1 0 x97 0 -1
Gyc1_98 y1 0 x98 0 -1
Gyc1_99 y1 0 x99 0 -1
Gyc1_100 y1 0 x100 0 -1
Gyc1_101 y1 0 x101 0 -1
Gyc1_102 y1 0 x102 0 -1
Gyc1_103 y1 0 x103 0 -1
Gyc1_104 y1 0 x104 0 -1
Gyc1_105 y1 0 x105 0 1
Gyc1_106 y1 0 x106 0 -1
Gyc1_107 y1 0 x107 0 1
Gyc1_108 y1 0 x108 0 -1
Gyc1_109 y1 0 x109 0 -1
Gyc1_110 y1 0 x110 0 -1
Gyc1_111 y1 0 x111 0 1
Gyc1_112 y1 0 x112 0 -1
Gyc1_113 y1 0 x113 0 1
Gyc1_114 y1 0 x114 0 -1
Gyc1_115 y1 0 x115 0 1
Gyc1_116 y1 0 x116 0 1
Gyc1_117 y1 0 x117 0 1
Gyc1_118 y1 0 x118 0 1
Gyc1_119 y1 0 x119 0 1
Gyc1_120 y1 0 x120 0 1
Gyc1_121 y1 0 x121 0 -1
Gyc1_122 y1 0 x122 0 -1
Gyc1_123 y1 0 x123 0 -1
Gyc1_124 y1 0 x124 0 1
Gyc1_125 y1 0 x125 0 -1
Gyc1_126 y1 0 x126 0 -1
Gyc1_127 y1 0 x127 0 -1
Gyc1_128 y1 0 x128 0 -1
Gyc1_129 y1 0 x129 0 -1
Gyc1_130 y1 0 x130 0 1
Gyc1_131 y1 0 x131 0 1
Gyc1_132 y1 0 x132 0 1
Gyc1_133 y1 0 x133 0 1
Gyc1_134 y1 0 x134 0 -1
Gyc1_135 y1 0 x135 0 -1
Gyc1_136 y1 0 x136 0 -1
Gyc1_137 y1 0 x137 0 1
Gyc1_138 y1 0 x138 0 -1
Gyc1_139 y1 0 x139 0 1
Gyc1_140 y1 0 x140 0 1
Gyc1_141 y1 0 x141 0 -1
Gyc1_142 y1 0 x142 0 -1
Gyc1_143 y1 0 x143 0 -1
Gyc1_144 y1 0 x144 0 1
Gyc1_145 y1 0 x145 0 1
Gyc1_146 y1 0 x146 0 1
Gyc1_147 y1 0 x147 0 0.640793612069572
Gyc1_148 y1 0 x148 0 -1
Gyc1_149 y1 0 x149 0 -1
Gyc1_150 y1 0 x150 0 -1
Gyc1_151 y1 0 x151 0 -1
Gyc1_152 y1 0 x152 0 1
Gyc1_153 y1 0 x153 0 -1
Gyc1_154 y1 0 x154 0 1
Gyc1_155 y1 0 x155 0 1
Gyc1_156 y1 0 x156 0 1
Gyc1_157 y1 0 x157 0 1
Gyc1_158 y1 0 x158 0 -1
Gyc1_159 y1 0 x159 0 1
Gyc1_160 y1 0 x160 0 0.507923162940901
Gyc1_161 y1 0 x161 0 -1
Gyc1_162 y1 0 x162 0 1
Gyc1_163 y1 0 x163 0 -1
Gyc1_164 y1 0 x164 0 -1
Gyc1_165 y1 0 x165 0 -1
Gyc1_166 y1 0 x166 0 -1
Gyc1_167 y1 0 x167 0 1
Gyc1_168 y1 0 x168 0 1
Gyc1_169 y1 0 x169 0 1
Gyc1_170 y1 0 x170 0 -1
Gyc1_171 y1 0 x171 0 1
Gyc1_172 y1 0 x172 0 1
Gyc1_173 y1 0 x173 0 -1
Gyc1_174 y1 0 x174 0 -1
Gyc1_175 y1 0 x175 0 1
Gyc1_176 y1 0 x176 0 1
Gyc1_177 y1 0 x177 0 -1
Gyc1_178 y1 0 x178 0 1
Gyc1_179 y1 0 x179 0 1
Gyc1_180 y1 0 x180 0 -1
Gyc1_181 y1 0 x181 0 -1
Gyc1_182 y1 0 x182 0 -1
Gyc1_183 y1 0 x183 0 1
Gyc1_184 y1 0 x184 0 -1
Gyc1_185 y1 0 x185 0 1
Gyc1_186 y1 0 x186 0 -1
Gyc1_187 y1 0 x187 0 -1
Gyc1_188 y1 0 x188 0 -1
Gyc1_189 y1 0 x189 0 -1
Gyc1_190 y1 0 x190 0 -1
Gyc1_191 y1 0 x191 0 -1
Gyc1_192 y1 0 x192 0 -1
Gyc1_193 y1 0 x193 0 1
Gyc1_194 y1 0 x194 0 1
Gyc1_195 y1 0 x195 0 1
Gyc1_196 y1 0 x196 0 -1
Gyc1_197 y1 0 x197 0 -1
Gyc1_198 y1 0 x198 0 1
Gyc1_199 y1 0 x199 0 -1
Gyc1_200 y1 0 x200 0 1
Gyc1_201 y1 0 x201 0 1
Gyc1_202 y1 0 x202 0 1
Gyc1_203 y1 0 x203 0 -1
Gyc1_204 y1 0 x204 0 1
Gyc1_205 y1 0 x205 0 -1
Gyc1_206 y1 0 x206 0 -1
Gyc1_207 y1 0 x207 0 1
Gyc1_208 y1 0 x208 0 1
Gyc1_209 y1 0 x209 0 -1
Gyc1_210 y1 0 x210 0 -1
Gyc1_211 y1 0 x211 0 -0.469538251234225
Gyc1_212 y1 0 x212 0 -1
Gyc1_213 y1 0 x213 0 -1
Gyc1_214 y1 0 x214 0 -1
Gyc1_215 y1 0 x215 0 -1
Gyc1_216 y1 0 x216 0 1
Gyc1_217 y1 0 x217 0 -1
Gyc1_218 y1 0 x218 0 -1
Gyc1_219 y1 0 x219 0 -1
Gyc1_220 y1 0 x220 0 1
Gyc1_221 y1 0 x221 0 1
Gyc1_222 y1 0 x222 0 -1
Gyc1_223 y1 0 x223 0 1
Gyc1_224 y1 0 x224 0 -1
Gyc1_225 y1 0 x225 0 -1
Gyc1_226 y1 0 x226 0 -1
Gyc1_227 y1 0 x227 0 1
Gyc1_228 y1 0 x228 0 -1
Gyc1_229 y1 0 x229 0 1
Gyc1_230 y1 0 x230 0 1
Gyc1_231 y1 0 x231 0 1
Gyc1_232 y1 0 x232 0 1
Gyc1_233 y1 0 x233 0 1
Gyc1_234 y1 0 x234 0 -1
Gyc1_235 y1 0 x235 0 -1
Gyc1_236 y1 0 x236 0 1
Gyc1_237 y1 0 x237 0 -1
Gyc1_238 y1 0 x238 0 1
Gyc1_239 y1 0 x239 0 -1
Gyc1_240 y1 0 x240 0 -1
Gyc1_241 y1 0 x241 0 -1
Gyc1_242 y1 0 x242 0 1
Gyc1_243 y1 0 x243 0 -1
Gyc1_244 y1 0 x244 0 1
Gyc1_245 y1 0 x245 0 -1
Gyc1_246 y1 0 x246 0 -1
Gyc1_247 y1 0 x247 0 1
Gyc1_248 y1 0 x248 0 1
Gyc1_249 y1 0 x249 0 -1
Gyc1_250 y1 0 x250 0 -1
Gyc1_251 y1 0 x251 0 1
Gyc1_252 y1 0 x252 0 1
Gyc1_253 y1 0 x253 0 -1
Gyc1_254 y1 0 x254 0 1
Gyc1_255 y1 0 x255 0 1
Gyc1_256 y1 0 x256 0 -1
Gyc1_257 y1 0 x257 0 -1
Gyc1_258 y1 0 x258 0 -1
Gyc1_259 y1 0 x259 0 1
Gyc1_260 y1 0 x260 0 -1
Gyc1_261 y1 0 x261 0 1
Gyc1_262 y1 0 x262 0 -1
Gyc1_263 y1 0 x263 0 1
Gyc1_264 y1 0 x264 0 -1
Gyc1_265 y1 0 x265 0 -1
Gyc1_266 y1 0 x266 0 -1
Gyc1_267 y1 0 x267 0 -1
Gyc1_268 y1 0 x268 0 1
Gyc1_269 y1 0 x269 0 1
Gyc1_270 y1 0 x270 0 1
Gyc1_271 y1 0 x271 0 1
Gyc1_272 y1 0 x272 0 -1
Gyc1_273 y1 0 x273 0 1
Gyc1_274 y1 0 x274 0 1
Gyc1_275 y1 0 x275 0 -1
Gyc1_276 y1 0 x276 0 1
Gyc1_277 y1 0 x277 0 -1
Gyc1_278 y1 0 x278 0 -1
Gyc1_279 y1 0 x279 0 1
Gyc1_280 y1 0 x280 0 1
Gyc1_281 y1 0 x281 0 1
Gyc1_282 y1 0 x282 0 -1
Gyc1_283 y1 0 x283 0 1
Gyc1_284 y1 0 x284 0 -1
Gyc1_285 y1 0 x285 0 1
Gyc1_286 y1 0 x286 0 -1
Gyc1_287 y1 0 x287 0 -1
Gyc1_288 y1 0 x288 0 1
Gyc1_289 y1 0 x289 0 -1
Gyc1_290 y1 0 x290 0 1
Gyc1_291 y1 0 x291 0 1
Gyc1_292 y1 0 x292 0 1
Gyc1_293 y1 0 x293 0 1
Gyc1_294 y1 0 x294 0 -1
Gyc1_295 y1 0 x295 0 -1
Gyc1_296 y1 0 x296 0 1
Gyc1_297 y1 0 x297 0 -1
Gyc1_298 y1 0 x298 0 1
Gyc1_299 y1 0 x299 0 -1
Gyc1_300 y1 0 x300 0 -1
Gyc1_301 y1 0 x301 0 -1
Gyc1_302 y1 0 x302 0 1
Gyc1_303 y1 0 x303 0 1
Gyc1_304 y1 0 x304 0 -1
Gyc1_305 y1 0 x305 0 1
Gyc1_306 y1 0 x306 0 1
Gyc1_307 y1 0 x307 0 1
Gyc1_308 y1 0 x308 0 -1
Gyc1_309 y1 0 x309 0 -1
Gyc1_310 y1 0 x310 0 -1
Gyc1_311 y1 0 x311 0 1
Gyc1_312 y1 0 x312 0 1
Gyc1_313 y1 0 x313 0 -0.520701327738653
Gyc1_314 y1 0 x314 0 1
Gyc1_315 y1 0 x315 0 1
Gyc1_316 y1 0 x316 0 1
Gyc1_317 y1 0 x317 0 -1
Gyc1_318 y1 0 x318 0 1
Gyc1_319 y1 0 x319 0 -1
Gyc1_320 y1 0 x320 0 1
Gyc1_321 y1 0 x321 0 1
Gyc1_322 y1 0 x322 0 1
Gyc1_323 y1 0 x323 0 -1
Gyc1_324 y1 0 x324 0 -1
Gyc1_325 y1 0 x325 0 -1
Gyc1_326 y1 0 x326 0 1
Gyc1_327 y1 0 x327 0 1
Gyc1_328 y1 0 x328 0 1
Gyc1_329 y1 0 x329 0 1
Gyc1_330 y1 0 x330 0 1
Gyc1_331 y1 0 x331 0 1
Gyc1_332 y1 0 x332 0 1
Gyc1_333 y1 0 x333 0 -1
Gyc1_334 y1 0 x334 0 1
Gyc1_335 y1 0 x335 0 1
Gyc1_336 y1 0 x336 0 1
Gyc1_337 y1 0 x337 0 1
Gyc1_338 y1 0 x338 0 1
Gyc1_339 y1 0 x339 0 -1
Gyc1_340 y1 0 x340 0 -1
Gyc1_341 y1 0 x341 0 1
Gyc1_342 y1 0 x342 0 1
Gyc1_343 y1 0 x343 0 1
Gyc1_344 y1 0 x344 0 1
Gyc1_345 y1 0 x345 0 1
Gyc1_346 y1 0 x346 0 -1
Gyc1_347 y1 0 x347 0 -1
Gyc1_348 y1 0 x348 0 1
Gyc1_349 y1 0 x349 0 1
Gyc1_350 y1 0 x350 0 1
Gyc1_351 y1 0 x351 0 -1
Gyc1_352 y1 0 x352 0 1
Gyc1_353 y1 0 x353 0 1
Gyc1_354 y1 0 x354 0 1
Gyc1_355 y1 0 x355 0 -1
Gyc1_356 y1 0 x356 0 -1
Gyc1_357 y1 0 x357 0 -1
Gyc1_358 y1 0 x358 0 -1
Gyc1_359 y1 0 x359 0 1
Gyc1_360 y1 0 x360 0 1
Gyc1_361 y1 0 x361 0 -0.0221922609234389
Gyc1_362 y1 0 x362 0 -1
Gyc1_363 y1 0 x363 0 -1
Gyc1_364 y1 0 x364 0 1
Gyc1_365 y1 0 x365 0 1
Gyc1_366 y1 0 x366 0 1
Gyc1_367 y1 0 x367 0 -1
Gyc1_368 y1 0 x368 0 -1
Gyc1_369 y1 0 x369 0 -1
Gyc1_370 y1 0 x370 0 -1
Gyc1_371 y1 0 x371 0 1
Gyc1_372 y1 0 x372 0 1
Gyc1_373 y1 0 x373 0 1
Gyc1_374 y1 0 x374 0 -0.384708635512887
Gyc1_375 y1 0 x375 0 1
Gyc1_376 y1 0 x376 0 -1
Gyc1_377 y1 0 x377 0 -1
Gyc1_378 y1 0 x378 0 1
Gyc1_379 y1 0 x379 0 -1
Gyc1_380 y1 0 x380 0 -1
Gyc1_381 y1 0 x381 0 -1
Gyc1_382 y1 0 x382 0 1
Gyc1_383 y1 0 x383 0 1
Gyc1_384 y1 0 x384 0 -1
Gyc1_385 y1 0 x385 0 -1
Gyc1_386 y1 0 x386 0 1
Gyc1_387 y1 0 x387 0 -1
Gyc1_388 y1 0 x388 0 1
Gyc1_389 y1 0 x389 0 -1
Gyc1_390 y1 0 x390 0 -1
Gyc1_391 y1 0 x391 0 1
Gyc1_392 y1 0 x392 0 -1
Gyc1_393 y1 0 x393 0 -1
Gyc1_394 y1 0 x394 0 -1
Gyc1_395 y1 0 x395 0 1
Gyc1_396 y1 0 x396 0 1
Gyc1_397 y1 0 x397 0 -1
Gyc1_398 y1 0 x398 0 -1
Gyc1_399 y1 0 x399 0 -1
Gyc1_400 y1 0 x400 0 1
Gyc1_401 y1 0 x401 0 1
Gyc1_402 y1 0 x402 0 -1
Gyc1_403 y1 0 x403 0 1
Gyc1_404 y1 0 x404 0 -1
Gyc1_405 y1 0 x405 0 1
Gyc1_406 y1 0 x406 0 1
Gyc1_407 y1 0 x407 0 -1
Gyc1_408 y1 0 x408 0 1
Gyc1_409 y1 0 x409 0 1
Gyc1_410 y1 0 x410 0 1
Gyc1_411 y1 0 x411 0 1
Gyc1_412 y1 0 x412 0 1
Gyc1_413 y1 0 x413 0 1
Gyc1_414 y1 0 x414 0 -1
Gyc1_415 y1 0 x415 0 1
Gyc1_416 y1 0 x416 0 1
Gyc1_417 y1 0 x417 0 -1
Gyc1_418 y1 0 x418 0 -1
Gyc1_419 y1 0 x419 0 -1
Gyc1_420 y1 0 x420 0 -1
Gyc1_421 y1 0 x421 0 1
Gyc1_422 y1 0 x422 0 -1
Gyc1_423 y1 0 x423 0 -0.744840083464683
Gyc1_424 y1 0 x424 0 -1
Gyc1_425 y1 0 x425 0 1
Gyc1_426 y1 0 x426 0 -1
Gyc1_427 y1 0 x427 0 1
Gyc1_428 y1 0 x428 0 -1
Gyc1_429 y1 0 x429 0 1
Gyc1_430 y1 0 x430 0 -1
Gyc1_431 y1 0 x431 0 -1
Gyc1_432 y1 0 x432 0 -1
Gyc1_433 y1 0 x433 0 1
Gyc1_434 y1 0 x434 0 -1
Gyc1_435 y1 0 x435 0 1
Gyc1_436 y1 0 x436 0 -1
Gyc1_437 y1 0 x437 0 -1
Gyc1_438 y1 0 x438 0 1
Gyc1_439 y1 0 x439 0 1
Gyc1_440 y1 0 x440 0 -1
Gyc1_441 y1 0 x441 0 1
Gyc1_442 y1 0 x442 0 1
Gyc1_443 y1 0 x443 0 -1
Gyc1_444 y1 0 x444 0 -1
Gyc1_445 y1 0 x445 0 -1
Gyc1_446 y1 0 x446 0 1
Gyc1_447 y1 0 x447 0 1
Gyc1_448 y1 0 x448 0 1
Gyc1_449 y1 0 x449 0 -1
Gyc1_450 y1 0 x450 0 1
Gyc1_451 y1 0 x451 0 1
Gyc1_452 y1 0 x452 0 1
Gyc1_453 y1 0 x453 0 -1
Gyc1_454 y1 0 x454 0 1
Gyc1_455 y1 0 x455 0 -1
Gyc1_456 y1 0 x456 0 -1
Gyc1_457 y1 0 x457 0 1
Gyc1_458 y1 0 x458 0 -1
Gyc1_459 y1 0 x459 0 -1
Gyc1_460 y1 0 x460 0 -1
Gyc1_461 y1 0 x461 0 1
Gyc1_462 y1 0 x462 0 -1
Gyc1_463 y1 0 x463 0 1
Gyc1_464 y1 0 x464 0 1
Gyc1_465 y1 0 x465 0 1
Gyc1_466 y1 0 x466 0 -1
Gyc1_467 y1 0 x467 0 1
Gyc1_468 y1 0 x468 0 1
Gyc1_469 y1 0 x469 0 -1
Gyc1_470 y1 0 x470 0 1
Gyc1_471 y1 0 x471 0 -1
Gyc1_472 y1 0 x472 0 -1
Gyc1_473 y1 0 x473 0 -1
Gyc1_474 y1 0 x474 0 -1
Gyc1_475 y1 0 x475 0 1
Gyc1_476 y1 0 x476 0 -1
Gyc1_477 y1 0 x477 0 1
Gyc1_478 y1 0 x478 0 -1
Gyc1_479 y1 0 x479 0 -1
Gyc1_480 y1 0 x480 0 -1
Gyc1_481 y1 0 x481 0 1
Gyc1_482 y1 0 x482 0 -1
Gyc1_483 y1 0 x483 0 1
Gyc1_484 y1 0 x484 0 1
Gyc1_485 y1 0 x485 0 1
Gyc1_486 y1 0 x486 0 1
Gyc1_487 y1 0 x487 0 -1
Gyc1_488 y1 0 x488 0 -1
Gyc1_489 y1 0 x489 0 1
Gyc1_490 y1 0 x490 0 -1
Gyc1_491 y1 0 x491 0 1
Gyc1_492 y1 0 x492 0 -1
Gyc1_493 y1 0 x493 0 1
Gyc1_494 y1 0 x494 0 1
Gyc1_495 y1 0 x495 0 1
Gyc1_496 y1 0 x496 0 1
Gyc1_497 y1 0 x497 0 -1
Gyc1_498 y1 0 x498 0 -1
Gyc1_499 y1 0 x499 0 -1
Gyc1_500 y1 0 x500 0 -1
Gyc1_501 y1 0 x501 0 1
Gyc1_502 y1 0 x502 0 -1
Gyc1_503 y1 0 x503 0 -1
Gyc1_504 y1 0 x504 0 -1
Gyc1_505 y1 0 x505 0 -1
Gyc1_506 y1 0 x506 0 1
Gyc1_507 y1 0 x507 0 1
Gyc1_508 y1 0 x508 0 1
Gyc1_509 y1 0 x509 0 1
Gyc1_510 y1 0 x510 0 1
Gyc1_511 y1 0 x511 0 -1
Gyc1_512 y1 0 x512 0 -1
Gyc1_513 y1 0 x513 0 1
Gyc1_514 y1 0 x514 0 -1
Gyc1_515 y1 0 x515 0 1
Gyc1_516 y1 0 x516 0 -1
Gyc1_517 y1 0 x517 0 -1
Gyc1_518 y1 0 x518 0 1
Gyc1_519 y1 0 x519 0 1
Gyc1_520 y1 0 x520 0 -1
Gyc1_521 y1 0 x521 0 1
Gyc1_522 y1 0 x522 0 -1
Gyc1_523 y1 0 x523 0 1
Gyc1_524 y1 0 x524 0 -1
Gyc1_525 y1 0 x525 0 1
Gyc1_526 y1 0 x526 0 -1
Gyc1_527 y1 0 x527 0 -1
Gyc1_528 y1 0 x528 0 1
Gyc1_529 y1 0 x529 0 1
Gyc1_530 y1 0 x530 0 -1
Gyc1_531 y1 0 x531 0 -1
Gyc1_532 y1 0 x532 0 1
Gyc1_533 y1 0 x533 0 1
Gyc1_534 y1 0 x534 0 -1
Gyc1_535 y1 0 x535 0 -1
Gyc1_536 y1 0 x536 0 1
Gyc1_537 y1 0 x537 0 1
Gyc1_538 y1 0 x538 0 1
Gyc1_539 y1 0 x539 0 1
Gyc1_540 y1 0 x540 0 1
Gyc1_541 y1 0 x541 0 -1
Gyc1_542 y1 0 x542 0 1
Gyc1_543 y1 0 x543 0 1
Gyc1_544 y1 0 x544 0 -1
Gyc1_545 y1 0 x545 0 1
Gyc1_546 y1 0 x546 0 -1
Gyc1_547 y1 0 x547 0 -1
Gyc1_548 y1 0 x548 0 -0.368747553746938
Gyc1_549 y1 0 x549 0 1
Gyc1_550 y1 0 x550 0 -1
Gyc1_551 y1 0 x551 0 1
Gyc1_552 y1 0 x552 0 -1
Gyc1_553 y1 0 x553 0 1
Gyc1_554 y1 0 x554 0 1
Gyc1_555 y1 0 x555 0 -1
Gyc1_556 y1 0 x556 0 -1
Gyc1_557 y1 0 x557 0 0.561328176894867
Gyc1_558 y1 0 x558 0 1
Gyc1_559 y1 0 x559 0 1
Gyc1_560 y1 0 x560 0 -1
Gyc1_561 y1 0 x561 0 -0.115207903522439
Gyc1_562 y1 0 x562 0 -1
Gyc1_563 y1 0 x563 0 1
Gyc1_564 y1 0 x564 0 -1
Gyc1_565 y1 0 x565 0 -1
Gyc1_566 y1 0 x566 0 1
Gyc1_567 y1 0 x567 0 -1
Gyc1_568 y1 0 x568 0 -1
Gyc1_569 y1 0 x569 0 -1
Gyc1_570 y1 0 x570 0 1
Gyc1_571 y1 0 x571 0 1
Gyc1_572 y1 0 x572 0 -1
Gyc1_573 y1 0 x573 0 1
Gyc1_574 y1 0 x574 0 1
Gyc1_575 y1 0 x575 0 -0.0994015716642623
Gyc1_576 y1 0 x576 0 1
Gyc1_577 y1 0 x577 0 1
Gyc1_578 y1 0 x578 0 -1
Gyc1_579 y1 0 x579 0 -1
Gyc1_580 y1 0 x580 0 1
Gyc1_581 y1 0 x581 0 1
Gyc1_582 y1 0 x582 0 -1
Gyc1_583 y1 0 x583 0 1
Gyc1_584 y1 0 x584 0 -1
Gyc1_585 y1 0 x585 0 1
Gyc1_586 y1 0 x586 0 -1
Gyc1_587 y1 0 x587 0 1
Gyc1_588 y1 0 x588 0 1
Gyc1_589 y1 0 x589 0 -1
Gyc1_590 y1 0 x590 0 -1
Gyc1_591 y1 0 x591 0 1
Gyc1_592 y1 0 x592 0 -1
Gyc1_593 y1 0 x593 0 -1
Gyc1_594 y1 0 x594 0 -1
Gyc1_595 y1 0 x595 0 -1
Gyc1_596 y1 0 x596 0 -1
Gyc1_597 y1 0 x597 0 1
Gyc1_598 y1 0 x598 0 -1
Gyc1_599 y1 0 x599 0 1
Gyc1_600 y1 0 x600 0 -1
Gyc1_601 y1 0 x601 0 -1
Gyc1_602 y1 0 x602 0 -1
Gyc1_603 y1 0 x603 0 -1
Gyc1_604 y1 0 x604 0 1
Gyc1_605 y1 0 x605 0 1
Gyc1_606 y1 0 x606 0 -1
Gyc1_607 y1 0 x607 0 1
Gyc1_608 y1 0 x608 0 1
Gyc1_609 y1 0 x609 0 1
Gyc1_610 y1 0 x610 0 1
Gyc1_611 y1 0 x611 0 -1
Gyc1_612 y1 0 x612 0 -1
Gyc1_613 y1 0 x613 0 -1
Gyc1_614 y1 0 x614 0 1
Gyc1_615 y1 0 x615 0 -1
Gyc1_616 y1 0 x616 0 -1
Gyc1_617 y1 0 x617 0 -1
Gyc1_618 y1 0 x618 0 1
Gyc1_619 y1 0 x619 0 -1
Gyc1_620 y1 0 x620 0 1
Gyc1_621 y1 0 x621 0 -1
Gyc1_622 y1 0 x622 0 1
Gyc1_623 y1 0 x623 0 1
Gyc1_624 y1 0 x624 0 -1
Gyc1_625 y1 0 x625 0 -1
Gyc1_626 y1 0 x626 0 -1
Gyc1_627 y1 0 x627 0 -1
Gyc1_628 y1 0 x628 0 1
Gyc1_629 y1 0 x629 0 1
Gyc1_630 y1 0 x630 0 1
Gyc1_631 y1 0 x631 0 1
Gyc1_632 y1 0 x632 0 -1
Gyc1_633 y1 0 x633 0 1
Gyc1_634 y1 0 x634 0 1
Gyc1_635 y1 0 x635 0 -1
Gyc1_636 y1 0 x636 0 -1
Gyc1_637 y1 0 x637 0 1
Gyc1_638 y1 0 x638 0 -1
Gyc1_639 y1 0 x639 0 -1
Gyc1_640 y1 0 x640 0 -1
Gyc1_641 y1 0 x641 0 -1
Gyc1_642 y1 0 x642 0 1
Gyc1_643 y1 0 x643 0 -1
Gyc1_644 y1 0 x644 0 1
Gyc1_645 y1 0 x645 0 -1
Gyc1_646 y1 0 x646 0 -1
Gyc1_647 y1 0 x647 0 -1
Gyc1_648 y1 0 x648 0 -1
Gyc1_649 y1 0 x649 0 1
Gyc1_650 y1 0 x650 0 -1
Gyc1_651 y1 0 x651 0 -1
Gyc1_652 y1 0 x652 0 -1
Gyc1_653 y1 0 x653 0 -1
Gyc1_654 y1 0 x654 0 -1
Gyc1_655 y1 0 x655 0 1
Gyc1_656 y1 0 x656 0 1
Gyc1_657 y1 0 x657 0 -1
Gyc1_658 y1 0 x658 0 -1
Gyc1_659 y1 0 x659 0 1
Gyc1_660 y1 0 x660 0 1
Gyc1_661 y1 0 x661 0 1
Gyc1_662 y1 0 x662 0 1
Gyc1_663 y1 0 x663 0 -1
Gyc1_664 y1 0 x664 0 -1
Gyc1_665 y1 0 x665 0 1
Gyc1_666 y1 0 x666 0 1
Gyc1_667 y1 0 x667 0 -1
Gyc1_668 y1 0 x668 0 1
Gyc1_669 y1 0 x669 0 -1
Gyc1_670 y1 0 x670 0 -1
Gyc1_671 y1 0 x671 0 -1
Gyc1_672 y1 0 x672 0 1
Gyc1_673 y1 0 x673 0 -1
Gyc1_674 y1 0 x674 0 -1
Gyc1_675 y1 0 x675 0 1
Gyc1_676 y1 0 x676 0 1
Gyc1_677 y1 0 x677 0 1
Gyc1_678 y1 0 x678 0 -1
Gyc1_679 y1 0 x679 0 1
Gyc1_680 y1 0 x680 0 -1
Gyc1_681 y1 0 x681 0 1
Gyc1_682 y1 0 x682 0 1
Gyc1_683 y1 0 x683 0 -1
Gyc1_684 y1 0 x684 0 1
Gyc1_685 y1 0 x685 0 1
Gyc1_686 y1 0 x686 0 1
Gyc1_687 y1 0 x687 0 1
Gyc1_688 y1 0 x688 0 1
Gyc1_689 y1 0 x689 0 1
Gyc1_690 y1 0 x690 0 -0.429651368108745
Gyc1_691 y1 0 x691 0 1
Gyc1_692 y1 0 x692 0 1
Gyc1_693 y1 0 x693 0 1
Gyc1_694 y1 0 x694 0 -1
Gyc1_695 y1 0 x695 0 -1
Gyc1_696 y1 0 x696 0 -1
Gyc1_697 y1 0 x697 0 -1
Gyc1_698 y1 0 x698 0 -1
Gyc1_699 y1 0 x699 0 -0.0880374124173457
Gyc1_700 y1 0 x700 0 1
Gyc1_701 y1 0 x701 0 1
Gyc1_702 y1 0 x702 0 -1
Gyc1_703 y1 0 x703 0 -1
Gyc1_704 y1 0 x704 0 -1
Gyc1_705 y1 0 x705 0 -1
Gyc1_706 y1 0 x706 0 1
Gyc1_707 y1 0 x707 0 -1
Gyc1_708 y1 0 x708 0 1
Gyc1_709 y1 0 x709 0 -1
Gyc1_710 y1 0 x710 0 1
Gyc1_711 y1 0 x711 0 1
Gyc1_712 y1 0 x712 0 -1
Gyc1_713 y1 0 x713 0 -1
Gyc1_714 y1 0 x714 0 0.739300995024409
Gyc1_715 y1 0 x715 0 -1
Gyc1_716 y1 0 x716 0 1
Gyc1_717 y1 0 x717 0 1
Gyc1_718 y1 0 x718 0 -1
Gyc1_719 y1 0 x719 0 -1
Gyc1_720 y1 0 x720 0 -1
Gyc1_721 y1 0 x721 0 1
Gyc1_722 y1 0 x722 0 1
Gyc1_723 y1 0 x723 0 -1
Gyc1_724 y1 0 x724 0 -1
Gyc1_725 y1 0 x725 0 -1
Gyc1_726 y1 0 x726 0 1
Gyc1_727 y1 0 x727 0 1
Gyc1_728 y1 0 x728 0 -1
Gyc1_729 y1 0 x729 0 -1
Gyc1_730 y1 0 x730 0 1
Gyc1_731 y1 0 x731 0 -1
Gyc1_732 y1 0 x732 0 1
Gyc1_733 y1 0 x733 0 1
Gyc1_734 y1 0 x734 0 1
Gyc1_735 y1 0 x735 0 0.44626266192832
Gyc1_736 y1 0 x736 0 -1
Gyc1_737 y1 0 x737 0 1
Gyc1_738 y1 0 x738 0 1
Gyc1_739 y1 0 x739 0 1
Gyc1_740 y1 0 x740 0 1
Gyc1_741 y1 0 x741 0 1
Gyc1_742 y1 0 x742 0 -1
Gyc1_743 y1 0 x743 0 1
Gyc1_744 y1 0 x744 0 1
Gyc1_745 y1 0 x745 0 -1
Gyc1_746 y1 0 x746 0 -1
Gyc1_747 y1 0 x747 0 -1
Gyc1_748 y1 0 x748 0 -0.129342348742683
Gyc1_749 y1 0 x749 0 -1
Gyc1_750 y1 0 x750 0 1
Gyc1_751 y1 0 x751 0 -1
Gyc1_752 y1 0 x752 0 -1
Gyc1_753 y1 0 x753 0 -1
Gyc1_754 y1 0 x754 0 1
Gyc1_755 y1 0 x755 0 1
Gyc1_756 y1 0 x756 0 -1
Gyc1_757 y1 0 x757 0 1
Gyc1_758 y1 0 x758 0 1
Gyc1_759 y1 0 x759 0 1
Gyc1_760 y1 0 x760 0 -1
Gyc1_761 y1 0 x761 0 1
Gyc1_762 y1 0 x762 0 -1
Gyc1_763 y1 0 x763 0 -1
Gyc1_764 y1 0 x764 0 -1
Gyc1_765 y1 0 x765 0 1
Gyc1_766 y1 0 x766 0 1
Gyc1_767 y1 0 x767 0 -1
Gyc1_768 y1 0 x768 0 1
Gyc1_769 y1 0 x769 0 1
Gyc1_770 y1 0 x770 0 -1
Gyc1_771 y1 0 x771 0 1
Gyc1_772 y1 0 x772 0 1
Gyc1_773 y1 0 x773 0 1
Gyc1_774 y1 0 x774 0 1
Gyc1_775 y1 0 x775 0 1
Gyc1_776 y1 0 x776 0 1
Gyc1_777 y1 0 x777 0 -1
Gyc1_778 y1 0 x778 0 1
Gyc1_779 y1 0 x779 0 1
Gyc1_780 y1 0 x780 0 -1
Gyc1_781 y1 0 x781 0 1
Gyc1_782 y1 0 x782 0 1
Gyc1_783 y1 0 x783 0 1
Gyc1_784 y1 0 x784 0 -1
Gyc1_785 y1 0 x785 0 1
Gyc1_786 y1 0 x786 0 -1
Gyc1_787 y1 0 x787 0 -1
Gyc1_788 y1 0 x788 0 -1
Gyc1_789 y1 0 x789 0 -1
Gyc1_790 y1 0 x790 0 -1
Gyc1_791 y1 0 x791 0 -1
Gyc1_792 y1 0 x792 0 -1
Gyc1_793 y1 0 x793 0 -1
Gyc1_794 y1 0 x794 0 1
Gyc1_795 y1 0 x795 0 -1
Gyc1_796 y1 0 x796 0 -1
Gyc1_797 y1 0 x797 0 1
Gyc1_798 y1 0 x798 0 1
Gyc1_799 y1 0 x799 0 -1
Gyc1_800 y1 0 x800 0 1
Gyc1_801 y1 0 x801 0 -1
Gyc1_802 y1 0 x802 0 -0.0184985327953721
Gyc1_803 y1 0 x803 0 0.0184110629126407
Gyc1_804 y1 0 x804 0 -0.0162436821571664
Gyc1_805 y1 0 x805 0 -0.0306045996268399
Gyc1_806 y1 0 x806 0 -0.0185373915017361
Gyc1_807 y1 0 x807 0 0.189070072062709
Gyc1_808 y1 0 x808 0 0.0414733080274735
Gyc1_809 y1 0 x809 0 -0.0215762453612865
Gyc1_810 y1 0 x810 0 0.0327547369549518
Gyc1_811 y1 0 x811 0 0.102266230076766
Gyc1_812 y1 0 x812 0 0.0396111877104231
Gyc1_813 y1 0 x813 0 0.0182248418193239
Gyc1_814 y1 0 x814 0 -0.0426652333041768
Gyc1_815 y1 0 x815 0 0.0233307672914821
Gyc1_816 y1 0 x816 0 -0.0254223121664125
Gyc1_817 y1 0 x817 0 0.0317026848158787
Gyc1_818 y1 0 x818 0 -0.0422341979490574
Gyc1_819 y1 0 x819 0 -0.865340283181575
Gyc1_820 y1 0 x820 0 0.0206001035174261
Gyc1_821 y1 0 x821 0 0.0332907524162984
Gyc1_822 y1 0 x822 0 -0.0202246343274757
Gyc1_823 y1 0 x823 0 -0.0449365142456012
Gyc1_824 y1 0 x824 0 -0.0319421491999584
Gyc1_825 y1 0 x825 0 -0.0773056440293557
Gyc1_826 y1 0 x826 0 -0.0366205741610145
Gyc1_827 y1 0 x827 0 0.0229625533241089
Gyc1_828 y1 0 x828 0 -0.0665546380953982
Gyc1_829 y1 0 x829 0 0.025336330342546
Gyc1_830 y1 0 x830 0 -0.0357773659450906
Gyc1_831 y1 0 x831 0 0.0191362736612837
Gyc1_832 y1 0 x832 0 -0.0377955084794261
Gyc1_833 y1 0 x833 0 0.0212196971563052
Gyc1_834 y1 0 x834 0 -0.0331606236220865
Gyc1_835 y1 0 x835 0 -0.0111544211357252
Gyc1_836 y1 0 x836 0 0.0140293170221055
Gyc1_837 y1 0 x837 0 -0.0325183179966366
Gyc1_838 y1 0 x838 0 0.0284472231556788
Gyc1_839 y1 0 x839 0 -0.00854764331161664
Gyc1_840 y1 0 x840 0 0.0275110760289382
Gyc1_841 y1 0 x841 0 0.0599599595230354
Gyc1_842 y1 0 x842 0 -0.0381802179503219
Gyc1_843 y1 0 x843 0 0.0242465767683883
Gyc1_844 y1 0 x844 0 -0.0441561237813757
Gyc1_845 y1 0 x845 0 0.0490184931859496
Gyc1_846 y1 0 x846 0 -0.0337260025012186
Gyc1_847 y1 0 x847 0 -0.101036094834031
Gyc1_848 y1 0 x848 0 -0.0351407850802222
Gyc1_849 y1 0 x849 0 -0.0567537346538817
Gyc1_850 y1 0 x850 0 -0.0532750101998565
Gyc1_851 y1 0 x851 0 0.0456654314401564
Gyc1_852 y1 0 x852 0 0.0273393152842214
Gyc1_853 y1 0 x853 0 0.0339740653495366
Gyc1_854 y1 0 x854 0 -0.0304602935183633
Gyc1_855 y1 0 x855 0 0.0355927562300585
Gyc1_856 y1 0 x856 0 -0.0293050022707103
Gyc1_857 y1 0 x857 0 -0.0183799311108693
Gyc1_858 y1 0 x858 0 0.0319902745556987
Gyc1_859 y1 0 x859 0 -0.0111274297524853
Gyc1_860 y1 0 x860 0 -0.0211209641478713
Gyc1_861 y1 0 x861 0 -0.0316214615781104
Gyc1_862 y1 0 x862 0 0.0392700708831647
Gyc1_863 y1 0 x863 0 -0.10391266403583
Gyc1_864 y1 0 x864 0 0.00104918500141694
Gyc1_865 y1 0 x865 0 0.02358917440259
Gyc1_866 y1 0 x866 0 0.00332747037417315
Gyc1_867 y1 0 x867 0 0.0271610742657155
Gyc1_868 y1 0 x868 0 -0.0673029742984706
Gyc1_869 y1 0 x869 0 -0.00299233791088585
Gyc1_870 y1 0 x870 0 -0.034676969229843
Gyc1_871 y1 0 x871 0 -0.0384175175938943
Gyc1_872 y1 0 x872 0 -0.00905358989463042
Gyc1_873 y1 0 x873 0 -0.042338979792386
Gyc1_874 y1 0 x874 0 0.0207983337091121
Gyc1_875 y1 0 x875 0 -0.0590022158354968
Gyc1_876 y1 0 x876 0 -0.00858475982476788
Gyc1_877 y1 0 x877 0 -0.0324034507792318
Gyc1_878 y1 0 x878 0 0.0211960075184822
Gyc1_879 y1 0 x879 0 0.0177001650583581
Gyc1_880 y1 0 x880 0 -0.0196702430839494
Gyc1_881 y1 0 x881 0 0.0230136794296102
Gyc1_882 y1 0 x882 0 -0.00504981793743012
Gyc1_883 y1 0 x883 0 -0.0103819134387604
Gyc1_884 y1 0 x884 0 -0.0322771386842084
Gyc1_885 y1 0 x885 0 -0.62031215078925
Gyc1_886 y1 0 x886 0 0.0211634786107699
Gyc1_887 y1 0 x887 0 0.0207118695492898
Gyc1_888 y1 0 x888 0 0.493817633528618
Gyc1_889 y1 0 x889 0 -0.16198333359946
Gyc1_890 y1 0 x890 0 0.0716333361304253
Gyc1_891 y1 0 x891 0 0.0307418007729381
Gyc1_892 y1 0 x892 0 0.0282853209494329
Gyc1_893 y1 0 x893 0 1
Gyc1_894 y1 0 x894 0 0.0535800496169478
Gyc1_895 y1 0 x895 0 -0.0216634919343863
Gyc1_896 y1 0 x896 0 -0.032775469865282
Gyc1_897 y1 0 x897 0 -0.0241706099574562
Gyc1_898 y1 0 x898 0 -0.0134562188320602
Gyc1_899 y1 0 x899 0 -0.0304115174914069
Gyc1_900 y1 0 x900 0 -0.0396610230584437
Gyc1_901 y1 0 x901 0 -1
Gyc1_902 y1 0 x902 0 -0.0199454620344677
Gyc1_903 y1 0 x903 0 -0.0418450649136348
Gyc1_904 y1 0 x904 0 -0.0113738414032618
Gyc1_905 y1 0 x905 0 -0.0353902380598805
Gyc1_906 y1 0 x906 0 0.0315178727610856
Gyc1_907 y1 0 x907 0 -0.0137728423312669
Gyc1_908 y1 0 x908 0 0.0350305135609045
Gyc1_909 y1 0 x909 0 -0.00454900258104212
Gyc1_910 y1 0 x910 0 -0.0104080553733159
Gyc1_911 y1 0 x911 0 -0.0734602442426313
Gyc1_912 y1 0 x912 0 0.0190472442617414
Gyc1_913 y1 0 x913 0 -0.0231352383976961
Gyc1_914 y1 0 x914 0 0.0260524461187888
Gyc1_915 y1 0 x915 0 -0.0290712409091076
Gyc1_916 y1 0 x916 0 0.0767337705511673
Gyc1_917 y1 0 x917 0 0.0285219038244124
Gyc1_918 y1 0 x918 0 0.0200325776762134
Gyc1_919 y1 0 x919 0 0.0264082259285396
Gyc1_920 y1 0 x920 0 0.0272116236548483
Gyc1_921 y1 0 x921 0 0.0247137079415455
Gyc1_922 y1 0 x922 0 -0.0451042386013274
Gyc1_923 y1 0 x923 0 -0.0303169279739388
Gyc1_924 y1 0 x924 0 -0.0560153806796329
Gyc1_925 y1 0 x925 0 0.054176957768437
Gyc1_926 y1 0 x926 0 -0.0284648187591079
Gyc1_927 y1 0 x927 0 -0.0390048188644007
Gyc1_928 y1 0 x928 0 -0.0394911000948911
Gyc1_929 y1 0 x929 0 -0.0355096713077262
Gyc1_930 y1 0 x930 0 -0.0331490412542296
Gyc1_931 y1 0 x931 0 0.100815007847331
Gyc1_932 y1 0 x932 0 -0.0515269546531856
Gyc1_933 y1 0 x933 0 0.0586758914788004
Gyc1_934 y1 0 x934 0 0.0285768065157269
Gyc1_935 y1 0 x935 0 -0.0217772845425289
Gyc1_936 y1 0 x936 0 -0.0299597442735522
Gyc1_937 y1 0 x937 0 -0.0329544760398509
Gyc1_938 y1 0 x938 0 0.0256234338554223
Gyc1_939 y1 0 x939 0 -0.0275157196834185
Gyc1_940 y1 0 x940 0 0.0170720366492818
Gyc1_941 y1 0 x941 0 0.0145562195333909
Gyc1_942 y1 0 x942 0 -0.0282756507618615
Gyc1_943 y1 0 x943 0 -0.0353872315583598
Gyc1_944 y1 0 x944 0 -0.0362412203522314
Gyc1_945 y1 0 x945 0 0.0168938993336012
Gyc1_946 y1 0 x946 0 0.0226852889796007
Gyc1_947 y1 0 x947 0 0.045870824316278
Gyc1_948 y1 0 x948 0 0.0824843881986445
Gyc1_949 y1 0 x949 0 -0.352818546970026
Gyc1_950 y1 0 x950 0 -0.0292094773326753
Gyc1_951 y1 0 x951 0 -0.116777778918874
Gyc1_952 y1 0 x952 0 -0.0336985632506323
Gyc1_953 y1 0 x953 0 0.0126771754074428
Gyc1_954 y1 0 x954 0 -0.0337462955454545
Gyc1_955 y1 0 x955 0 0.00641976844601356
Gyc1_956 y1 0 x956 0 0.025438572377367
Gyc1_957 y1 0 x957 0 0.038121902993775
Gyc1_958 y1 0 x958 0 0.339153550578161
Gyc1_959 y1 0 x959 0 -0.112784098644399
Gyc1_960 y1 0 x960 0 0.0282822694354439
Gyc1_961 y1 0 x961 0 -0.00730347354240904
Gyc1_962 y1 0 x962 0 -0.0544324814373458
Gyc1_963 y1 0 x963 0 0.0286323503989267
Gyc1_964 y1 0 x964 0 -0.0269112428170093
Gyc1_965 y1 0 x965 0 -0.030009484818426
Gyc1_966 y1 0 x966 0 -0.00156623514418963
Gyc1_967 y1 0 x967 0 -0.0993587864098731
Gyc1_968 y1 0 x968 0 -0.0754512429200196
Gyc1_969 y1 0 x969 0 0.0287204274782699
Gyc1_970 y1 0 x970 0 0.017224536881483
Gyc1_971 y1 0 x971 0 -0.0291762916421159
Gyc1_972 y1 0 x972 0 0.0308772759394462
Gyc1_973 y1 0 x973 0 0.0412456599739009
Gyc1_974 y1 0 x974 0 -0.0190735850423843
Gyc1_975 y1 0 x975 0 0.0127184086363897
Gyc1_976 y1 0 x976 0 0.025605188773503
Gyc1_977 y1 0 x977 0 0.0277208452453148
Gyc1_978 y1 0 x978 0 -0.0407779020702821
Gyc1_979 y1 0 x979 0 0.0217201416500759
Gyc1_980 y1 0 x980 0 0.024359742157628
Gyc1_981 y1 0 x981 0 -0.0319032324321506
Gyc1_982 y1 0 x982 0 -0.122205447957412
Gyc1_983 y1 0 x983 0 -0.00600238845689024
Gyc1_984 y1 0 x984 0 0.0160832691149045
Gyc1_985 y1 0 x985 0 -0.0319361479926495
Gyc1_986 y1 0 x986 0 0.0219093873067092
Gyc1_987 y1 0 x987 0 -0.0244904850987887
Gyc1_988 y1 0 x988 0 -0.0268896607899563
Gyc1_989 y1 0 x989 0 -0.0316530955433984
Gyc1_990 y1 0 x990 0 -0.0273972387610521
Gyc1_991 y1 0 x991 0 -0.0306365255554227
Gyc1_992 y1 0 x992 0 -0.0246051473776224
Gyc1_993 y1 0 x993 0 -0.0278089665246527
Gyc1_994 y1 0 x994 0 0.0271031204559595
Gyc1_995 y1 0 x995 0 0.0289403906283485
Gyc1_996 y1 0 x996 0 0.0347355081479142
Gyc1_997 y1 0 x997 0 -0.0369461558637051
Gyc1_998 y1 0 x998 0 -0.0194523510895639
Gyc1_999 y1 0 x999 0 0.347626205692782
Gyc1_1000 y1 0 x1000 0 -0.0244467773916046
Gyc1_1001 y1 0 x1001 0 0.0120048556673994
Gyc1_1002 y1 0 x1002 0 0.138198574630681
Gyc1_1003 y1 0 x1003 0 0.0354828720373891
Gyc1_1004 y1 0 x1004 0 -0.0296281779247966
Gyc1_1005 y1 0 x1005 0 0.0166862106296218
Gyc1_1006 y1 0 x1006 0 -0.0247549959209378
Gyc1_1007 y1 0 x1007 0 -0.00620265568942191
Gyc1_1008 y1 0 x1008 0 0.0285025886320004
Gyc1_1009 y1 0 x1009 0 -0.0274285883739891
Gyc1_1010 y1 0 x1010 0 -0.0219566398217244
Gyc1_1011 y1 0 x1011 0 -0.0261329280223452
Gyc1_1012 y1 0 x1012 0 -0.132143169050949
Gyc1_1013 y1 0 x1013 0 0.0817747417248397
Gyc1_1014 y1 0 x1014 0 -0.037829547364336
Gyc1_1015 y1 0 x1015 0 -0.0263944986322371
Gyc1_1016 y1 0 x1016 0 -0.0274922796810143
Gyc1_1017 y1 0 x1017 0 0.0257643275454355
Gyc1_1018 y1 0 x1018 0 -0.0275040964469227
Gyc1_1019 y1 0 x1019 0 -0.0245787287169711
Gyc1_1020 y1 0 x1020 0 -0.0250656840922994
Gyc1_1021 y1 0 x1021 0 0.0290858403175264
Gyc1_1022 y1 0 x1022 0 0.0343230850370314
Gyc1_1023 y1 0 x1023 0 -0.0207762080548217
Gyc1_1024 y1 0 x1024 0 -0.000820480212370323
Gyc1_1025 y1 0 x1025 0 -0.0240491549581153
Gyc1_1026 y1 0 x1026 0 0.020893320155285
Gyc1_1027 y1 0 x1027 0 0.0559844074518265
Gyc1_1028 y1 0 x1028 0 0.0162975850382673
Gyc1_1029 y1 0 x1029 0 -0.015575112133273
Gyc1_1030 y1 0 x1030 0 0.0559428134738894
Gyc1_1031 y1 0 x1031 0 -0.0335563311078887
Gyc1_1032 y1 0 x1032 0 -0.0157485554760179
Gyc1_1033 y1 0 x1033 0 0.0293072001476516
Gyc1_1034 y1 0 x1034 0 0.00190669823759585
Gyc1_1035 y1 0 x1035 0 0.0429360358494343
Gyc1_1036 y1 0 x1036 0 -0.0147756987140752
Gyc1_1037 y1 0 x1037 0 -0.0675454364190956
Gyc1_1038 y1 0 x1038 0 -0.0308748268777714
Gyc1_1039 y1 0 x1039 0 1
Gyc1_1040 y1 0 x1040 0 -0.04967963746973
Gyc1_1041 y1 0 x1041 0 -0.0415240447034286
Gyc1_1042 y1 0 x1042 0 -0.0364685811242365
Gyc1_1043 y1 0 x1043 0 0.0511829707141436
Gyc1_1044 y1 0 x1044 0 -0.0326637232780836
Gyc1_1045 y1 0 x1045 0 0.0830762655707478
Gyc1_1046 y1 0 x1046 0 0.0882374783243279
Gyc1_1047 y1 0 x1047 0 -0.00979108040700255
Gyc1_1048 y1 0 x1048 0 0.0893530261043168
Gyc1_1049 y1 0 x1049 0 0.0501345246284436
Gyc1_1050 y1 0 x1050 0 -0.0285711461510834
Gyc1_1051 y1 0 x1051 0 -0.02477548311055
Gyc1_1052 y1 0 x1052 0 0.0730314771765023
Gyc1_1053 y1 0 x1053 0 0.0345122851701485
Gyc1_1054 y1 0 x1054 0 -0.0182599665901559
Gyc1_1055 y1 0 x1055 0 0.0220745132670166
Gyc1_1056 y1 0 x1056 0 0.0195052786566659
Gyc1_1057 y1 0 x1057 0 -0.0343949337245629
Gyc1_1058 y1 0 x1058 0 -0.0390627080120133
Gyc1_1059 y1 0 x1059 0 -0.0258496784615005
Gyc1_1060 y1 0 x1060 0 0.0148068024970531
Gyc1_1061 y1 0 x1061 0 -0.0349132775057883
Gyc1_1062 y1 0 x1062 0 0.030972111774135
Gyc1_1063 y1 0 x1063 0 -0.186428237808215
Gyc1_1064 y1 0 x1064 0 -0.00414897206136495
Gyc1_1065 y1 0 x1065 0 -0.0285842857474428
Gyc1_1066 y1 0 x1066 0 -0.0273874316410241
Gyc1_1067 y1 0 x1067 0 0.00580746634204673
Gyc1_1068 y1 0 x1068 0 -0.000808833247785905
Gyc1_1069 y1 0 x1069 0 0.026636947357113
Gyc1_1070 y1 0 x1070 0 0.0132240312236573
Gyc1_1071 y1 0 x1071 0 0.0226793326183319
Gyc1_1072 y1 0 x1072 0 0.00977680921024747
Gyc1_1073 y1 0 x1073 0 -0.00064701488138197
Gyc1_1074 y1 0 x1074 0 0.256346037432277
Gyc1_1075 y1 0 x1075 0 0.0157941411654877
Gyc1_1076 y1 0 x1076 0 -0.00888542343800524
Gyc1_1077 y1 0 x1077 0 -0.0260461452769963
Gyc1_1078 y1 0 x1078 0 0.00356444690274648
Gyc1_1079 y1 0 x1079 0 -0.0197018149615921
Gyc1_1080 y1 0 x1080 0 0.321567197054508
Gyc1_1081 y1 0 x1081 0 -0.0046306825609244
Gyc1_1082 y1 0 x1082 0 0.0226217795142258
Gyc1_1083 y1 0 x1083 0 -0.0273847123910682
Gyc1_1084 y1 0 x1084 0 0.00248690933598018
Gyc1_1085 y1 0 x1085 0 -0.0305827046866981
Gyc1_1086 y1 0 x1086 0 0.0244722026433671
Gyc1_1087 y1 0 x1087 0 -0.0214835990789603
Gyc1_1088 y1 0 x1088 0 -0.0234860905368189
Gyc1_1089 y1 0 x1089 0 -0.00741509827110348
Gyc1_1090 y1 0 x1090 0 -0.00905141732079048
Gyc1_1091 y1 0 x1091 0 0.0349507984277899
Gyc1_1092 y1 0 x1092 0 0.0219865058547984
Gyc1_1093 y1 0 x1093 0 0.0231421891901114
Gyc1_1094 y1 0 x1094 0 0.0116861328156036
Gyc1_1095 y1 0 x1095 0 -0.117990128096692
Gyc1_1096 y1 0 x1096 0 -0.0144074175293483
Gyc1_1097 y1 0 x1097 0 0.0929021461721447
Gyc1_1098 y1 0 x1098 0 -0.0378360739270374
Gyc1_1099 y1 0 x1099 0 0.0230153244920915
Gyc1_1100 y1 0 x1100 0 -0.0160262391334373
Gyc1_1101 y1 0 x1101 0 -0.0200504362298308
Gyc1_1102 y1 0 x1102 0 -0.0015258235534791
Gyc1_1103 y1 0 x1103 0 -0.00606196148543281
Gyc1_1104 y1 0 x1104 0 0.0229457711434528
Gyc1_1105 y1 0 x1105 0 0.031712794751209
Gyc1_1106 y1 0 x1106 0 0.0215224960928338
Gyc1_1107 y1 0 x1107 0 0.0281966499123909
Gyc1_1108 y1 0 x1108 0 0.0260857530075692
Gyc1_1109 y1 0 x1109 0 0.018998976791381
Gyc1_1110 y1 0 x1110 0 -0.0210750465123269
Gyc1_1111 y1 0 x1111 0 -0.031504554985058
Gyc1_1112 y1 0 x1112 0 -0.049208630535884
Gyc1_1113 y1 0 x1113 0 0.020143580555018
Gyc1_1114 y1 0 x1114 0 -0.0532491735224948
Gyc1_1115 y1 0 x1115 0 0.0281687629207278
Gyc1_1116 y1 0 x1116 0 0.0167899989838125
Gyc1_1117 y1 0 x1117 0 0.0193811617182527
Gyc1_1118 y1 0 x1118 0 -0.0310515026933192
Gyc1_1119 y1 0 x1119 0 0.0383809355470936
Gyc1_1120 y1 0 x1120 0 -0.0333941541439189
Gyc1_1121 y1 0 x1121 0 0.0251120342308776
Gyc1_1122 y1 0 x1122 0 0.0264294122037744
Gyc1_1123 y1 0 x1123 0 0.0287907154397907
Gyc1_1124 y1 0 x1124 0 -0.00955025749291967
Gyc1_1125 y1 0 x1125 0 -0.0151982287332185
Gyc1_1126 y1 0 x1126 0 -0.0199634200987534
Gyc1_1127 y1 0 x1127 0 0.0504865843736375
Gyc1_1128 y1 0 x1128 0 0.0257632365031656
Gyc1_1129 y1 0 x1129 0 0.0244370957055262
Gyc1_1130 y1 0 x1130 0 0.0529074325250413
Gyc1_1131 y1 0 x1131 0 0.0178519370559603
Gyc1_1132 y1 0 x1132 0 0.0300851308845024
Gyc1_1133 y1 0 x1133 0 0.237152020112785
Gyc1_1134 y1 0 x1134 0 0.0024316072460511
Gyc1_1135 y1 0 x1135 0 0.306674548667915
Gyc1_1136 y1 0 x1136 0 0.0124072297315233
Gyc1_1137 y1 0 x1137 0 0.0205159445343591
Gyc1_1138 y1 0 x1138 0 -0.0083130662697612
Gyc1_1139 y1 0 x1139 0 -0.0123743543892008
Gyc1_1140 y1 0 x1140 0 0.0431155089522299
Gyc1_1141 y1 0 x1141 0 -0.0177530176263122
Gyc1_1142 y1 0 x1142 0 0.0100304646912864
Gyc1_1143 y1 0 x1143 0 -0.0471006218387666
Gyc1_1144 y1 0 x1144 0 0.0330419262239764
Gyc1_1145 y1 0 x1145 0 0.0190734373170231
Gyc1_1146 y1 0 x1146 0 0.0116927391212164
Gyc1_1147 y1 0 x1147 0 0.0188614434778869
Gyc1_1148 y1 0 x1148 0 -0.0193632497251981
Gyc1_1149 y1 0 x1149 0 0.024268153169993
Gyc1_1150 y1 0 x1150 0 0.0186115287058802
Gyc1_1151 y1 0 x1151 0 0.028393123452864
Gyc1_1152 y1 0 x1152 0 -0.0198226405767151
Gyc1_1153 y1 0 x1153 0 -0.0238276972512639
Gyc1_1154 y1 0 x1154 0 0.0215115390077716
Gyc1_1155 y1 0 x1155 0 0.0298060399843724
Gyc1_1156 y1 0 x1156 0 -0.00438018972963146
Gyc1_1157 y1 0 x1157 0 -0.0273797225539813
Gyc1_1158 y1 0 x1158 0 0.10613005603359
Gyc1_1159 y1 0 x1159 0 -0.0262745869447876
Gyc1_1160 y1 0 x1160 0 -0.0545838751806378
Gyc1_1161 y1 0 x1161 0 0.0118470947719147
Gyc1_1162 y1 0 x1162 0 -0.0211229652154852
Gyc1_1163 y1 0 x1163 0 -0.0580701812063002
Gyc1_1164 y1 0 x1164 0 -0.0332279845354004
Gyc1_1165 y1 0 x1165 0 0.0240946838924812
Gyc1_1166 y1 0 x1166 0 0.02487223068265
Gyc1_1167 y1 0 x1167 0 0.0302224094590469
Gyc1_1168 y1 0 x1168 0 -0.0324678566172625
Gyc1_1169 y1 0 x1169 0 -0.0437353698943204
Gyc1_1170 y1 0 x1170 0 -0.0358674492892006
Gyc1_1171 y1 0 x1171 0 -0.0300473998165971
Gyc1_1172 y1 0 x1172 0 0.0238007764231463
Gyc1_1173 y1 0 x1173 0 0.0271538323619072
Gyc1_1174 y1 0 x1174 0 0.0208495042208759
Gyc1_1175 y1 0 x1175 0 0.10679937809944
Gyc1_1176 y1 0 x1176 0 0.0204365600172786
Gyc1_1177 y1 0 x1177 0 -0.0466611200709841
Gyc1_1178 y1 0 x1178 0 -0.028807083182489
Gyc1_1179 y1 0 x1179 0 0.0240263778552013
Gyc1_1180 y1 0 x1180 0 -0.020026799780592
Gyc1_1181 y1 0 x1181 0 -0.049297404324707
Gyc1_1182 y1 0 x1182 0 0.103407313010965
Gyc1_1183 y1 0 x1183 0 0.0113889910812287
Gyc1_1184 y1 0 x1184 0 0.0299302635516084
Gyc1_1185 y1 0 x1185 0 -0.0247732129910957
Gyc1_1186 y1 0 x1186 0 -0.0295686406422275
Gyc1_1187 y1 0 x1187 0 0.0386650227809823
Gyc1_1188 y1 0 x1188 0 -0.0228325927745304
Gyc1_1189 y1 0 x1189 0 0.0467039946261285
Gyc1_1190 y1 0 x1190 0 0.010312295852589
Gyc1_1191 y1 0 x1191 0 -0.0308232936453738
Gyc1_1192 y1 0 x1192 0 0.00879962940379789
Gyc1_1193 y1 0 x1193 0 -0.0323841332882776
Gyc1_1194 y1 0 x1194 0 -0.0292856795632559
Gyc1_1195 y1 0 x1195 0 -0.0338612172906472
Gyc1_1196 y1 0 x1196 0 -0.026086512560574
Gyc1_1197 y1 0 x1197 0 0.0287485342151601
Gyc1_1198 y1 0 x1198 0 -0.0219699995876249
Gyc1_1199 y1 0 x1199 0 -0.0307702393633883
Gyc1_1200 y1 0 x1200 0 0.00261327730692243
Gyc1_1201 y1 0 x1201 0 0.0338822700145655
Gyc1_1202 y1 0 x1202 0 0.0294885291134203
Gyc1_1203 y1 0 x1203 0 -0.0139670392716263
Gyc1_1204 y1 0 x1204 0 0.0279835264404544
Gyc1_1205 y1 0 x1205 0 -0.00461186287031922
Gyc1_1206 y1 0 x1206 0 0.0508673698720286
Gyc1_1207 y1 0 x1207 0 0.0220757238497013
Gyc1_1208 y1 0 x1208 0 -0.0404995973983076
Gyc1_1209 y1 0 x1209 0 0.027941149789188
Gyc1_1210 y1 0 x1210 0 0.20180918706796
Gyc1_1211 y1 0 x1211 0 -0.00758781857179836
Gyc1_1212 y1 0 x1212 0 0.0137678691582264
Gyc1_1213 y1 0 x1213 0 0.0322191615568716
Gyc1_1214 y1 0 x1214 0 0.0426299850081161
Gyc1_1215 y1 0 x1215 0 -0.055108969634416
Gyc1_1216 y1 0 x1216 0 0.0193620844116145
Gyc1_1217 y1 0 x1217 0 0.029327569302809
Gyc1_1218 y1 0 x1218 0 -0.044401752606949
Gyc1_1219 y1 0 x1219 0 -0.0222978675936387
Gyc1_1220 y1 0 x1220 0 -0.0298134125781267
Gyc1_1221 y1 0 x1221 0 -0.0366499432344821
Gyc1_1222 y1 0 x1222 0 0.0253488608456527
Gyc1_1223 y1 0 x1223 0 -0.257705049683437
Gyc1_1224 y1 0 x1224 0 -0.0387215721818984
Gyc1_1225 y1 0 x1225 0 -0.070772560929037
Gyc1_1226 y1 0 x1226 0 0.0180365216723429
Gyc1_1227 y1 0 x1227 0 -0.0301808526321762
Gyc1_1228 y1 0 x1228 0 0.0154456119551467
Gyc1_1229 y1 0 x1229 0 -0.0329812002860578
Gyc1_1230 y1 0 x1230 0 0.0250472684533126
Gyc1_1231 y1 0 x1231 0 -0.0237910977957059
Gyc1_1232 y1 0 x1232 0 -0.0220754318195815
Gyc1_1233 y1 0 x1233 0 -0.016190058591059
Gyc1_1234 y1 0 x1234 0 0.0218367649606027
Gyc1_1235 y1 0 x1235 0 -0.0321856501293208
Gyc1_1236 y1 0 x1236 0 0.0230988710980261
Gyc1_1237 y1 0 x1237 0 -0.00902986352171001
Gyc1_1238 y1 0 x1238 0 -0.0174077855573478
Gyc1_1239 y1 0 x1239 0 0.0257079648307056
Gyc1_1240 y1 0 x1240 0 0.0152379648738294
Gyc1_1241 y1 0 x1241 0 -0.0492359199659982
Gyc1_1242 y1 0 x1242 0 0.0282011690200929
Gyc1_1243 y1 0 x1243 0 0.0225172452483065
Gyc1_1244 y1 0 x1244 0 -0.0220311036592284
Gyc1_1245 y1 0 x1245 0 -0.017600197614151
Gyc1_1246 y1 0 x1246 0 -0.00351882246671352
Gyc1_1247 y1 0 x1247 0 -0.0167023457038029
Gyc1_1248 y1 0 x1248 0 0.0219540599463292
Gyc1_1249 y1 0 x1249 0 0.025044763497549
Gyc1_1250 y1 0 x1250 0 -0.0257926330841533
Gyc1_1251 y1 0 x1251 0 0.0214570574353549
Gyc1_1252 y1 0 x1252 0 0.451323918002395
Gyc1_1253 y1 0 x1253 0 0.0146312105547419
Gyc1_1254 y1 0 x1254 0 -0.0228298200235836
Gyc1_1255 y1 0 x1255 0 0.0208914897059767
Gyc1_1256 y1 0 x1256 0 -0.0205505357382281
Gyc1_1257 y1 0 x1257 0 -0.0111075859419247
Gyc1_1258 y1 0 x1258 0 0.0219521713164051
Gyc1_1259 y1 0 x1259 0 -0.0221820419429071
Gyc1_1260 y1 0 x1260 0 -0.022200411336219
Gyc1_1261 y1 0 x1261 0 -0.0252640723195727
Gyc1_1262 y1 0 x1262 0 0.0132995815708065
Gyc1_1263 y1 0 x1263 0 0.0106091070124245
Gyc1_1264 y1 0 x1264 0 0.0154030936489154
Gyc1_1265 y1 0 x1265 0 0.0112337394092409
Gyc1_1266 y1 0 x1266 0 0.0101838179336324
Gyc1_1267 y1 0 x1267 0 -0.00888007277393451
Gyc1_1268 y1 0 x1268 0 -0.560284341289593
Gyc1_1269 y1 0 x1269 0 0.02847821827518
Gyc1_1270 y1 0 x1270 0 -0.0243273079724769
Gyc1_1271 y1 0 x1271 0 0.0195180839610911
Gyc1_1272 y1 0 x1272 0 -0.0141965731214775
Gyc1_1273 y1 0 x1273 0 -0.0255530821402425
Gyc1_1274 y1 0 x1274 0 0.0553385428201636
Gyc1_1275 y1 0 x1275 0 -0.0244514132752405
Gyc1_1276 y1 0 x1276 0 0.0141152535504384
Gyc1_1277 y1 0 x1277 0 -0.0179399205837868
Gyc1_1278 y1 0 x1278 0 0.0175487786665809
Gyc1_1279 y1 0 x1279 0 -0.0243244278282056
Gyc1_1280 y1 0 x1280 0 -0.0266951991179635
Gyc1_1281 y1 0 x1281 0 -0.0183726122755261
Gyc1_1282 y1 0 x1282 0 0.0534294475354203
Gyc1_1283 y1 0 x1283 0 -0.0174599850413483
Gyc1_1284 y1 0 x1284 0 0.0238964620613008
Gyc1_1285 y1 0 x1285 0 0.0383561370775833
Gyc1_1286 y1 0 x1286 0 -0.0527887367171682
Gyc1_1287 y1 0 x1287 0 -0.0215890887617336
Gyc1_1288 y1 0 x1288 0 -0.0293107528114341
Gyc1_1289 y1 0 x1289 0 -0.0299305273902352
Gyc1_1290 y1 0 x1290 0 0.0380247721728445
Gyc1_1291 y1 0 x1291 0 -0.0352230822329012
Gyc1_1292 y1 0 x1292 0 0.00177684308972818
Gyc1_1293 y1 0 x1293 0 0.0190728276689542
Gyc1_1294 y1 0 x1294 0 0.0332232721508427
Gyc1_1295 y1 0 x1295 0 0.0245828651190196
Gyc1_1296 y1 0 x1296 0 0.013576544186524
Gyc1_1297 y1 0 x1297 0 0.0145801164317319
Gyc1_1298 y1 0 x1298 0 -0.00631933406204309
Gyc1_1299 y1 0 x1299 0 -0.0246823675196354
Gyc1_1300 y1 0 x1300 0 -0.0253297631917343
Gyc1_1301 y1 0 x1301 0 -0.00893944519136534
Gyc1_1302 y1 0 x1302 0 -0.153485621873898
Gyc1_1303 y1 0 x1303 0 -0.196102760450646
Gyc1_1304 y1 0 x1304 0 -0.0177459186755715
Gyc1_1305 y1 0 x1305 0 -0.0889243752057754
Gyc1_1306 y1 0 x1306 0 -0.0223061602641286
Gyc1_1307 y1 0 x1307 0 0.00479704045986906
Gyc1_1308 y1 0 x1308 0 0.0862715897012198
Gyc1_1309 y1 0 x1309 0 0.0240407692575535
Gyc1_1310 y1 0 x1310 0 0.06085710447896
Gyc1_1311 y1 0 x1311 0 0.00732883920974459
Gyc1_1312 y1 0 x1312 0 -0.0262352562918183
Gyc1_1313 y1 0 x1313 0 -0.0294375939153124
Gyc1_1314 y1 0 x1314 0 0.0246455105374502
Gyc1_1315 y1 0 x1315 0 -0.0155970012166573
Gyc1_1316 y1 0 x1316 0 -0.14478293193291
Gyc1_1317 y1 0 x1317 0 -0.0124372692389488
Gyc1_1318 y1 0 x1318 0 -0.020462359590545
Gyc1_1319 y1 0 x1319 0 -0.0623281275525448
Gyc1_1320 y1 0 x1320 0 0.019495681835295
Gyc1_1321 y1 0 x1321 0 -0.0162048867387543
Gyc1_1322 y1 0 x1322 0 0.0605779317190687
Gyc1_1323 y1 0 x1323 0 -0.00829776649561237
Gyc1_1324 y1 0 x1324 0 0.0273467902504997
Gyc1_1325 y1 0 x1325 0 -0.00900644211360539
Gyc1_1326 y1 0 x1326 0 0.0232623333513451
Gyc1_1327 y1 0 x1327 0 -0.0257527543895146
Gyc1_1328 y1 0 x1328 0 -0.0259362573272841
Gyc1_1329 y1 0 x1329 0 -0.0842025535184021
Gyc1_1330 y1 0 x1330 0 0.0251668369520219
Gyc1_1331 y1 0 x1331 0 -0.0143147229650577
Gyc1_1332 y1 0 x1332 0 -0.0177932436385091
Gyc1_1333 y1 0 x1333 0 0.0311973752702724
Gyc1_1334 y1 0 x1334 0 0.0275756595246855
Gyc1_1335 y1 0 x1335 0 0.081148949986509
Gyc1_1336 y1 0 x1336 0 -0.0238496571554055
Gyc1_1337 y1 0 x1337 0 0.0399428065995687
Gyc1_1338 y1 0 x1338 0 -0.02261323579782
Gyc1_1339 y1 0 x1339 0 0.0339487605222749
Gyc1_1340 y1 0 x1340 0 -0.0287366371969011
Gyc1_1341 y1 0 x1341 0 -0.0256725259637402
Gyc1_1342 y1 0 x1342 0 -0.020369001664095
Gyc1_1343 y1 0 x1343 0 0.0248248027559589
Gyc1_1344 y1 0 x1344 0 0.0247650510322117
Gyc1_1345 y1 0 x1345 0 0.0673717162857146
Gyc1_1346 y1 0 x1346 0 -0.0362672732803287
Gyc1_1347 y1 0 x1347 0 -0.0252292608923669
Gyc1_1348 y1 0 x1348 0 0.00276738036458263
Gyc1_1349 y1 0 x1349 0 0.0916568887885562
Gyc1_1350 y1 0 x1350 0 0.0367242517253528
Gyc1_1351 y1 0 x1351 0 -0.0220240280601424
Gyc1_1352 y1 0 x1352 0 0.0458890728942886
Gyc1_1353 y1 0 x1353 0 -0.0152549429774666
Gyc1_1354 y1 0 x1354 0 0.0102252964236384
Gyc1_1355 y1 0 x1355 0 0.0278454055908607
Gyc1_1356 y1 0 x1356 0 -0.00606615531396618
Gyc1_1357 y1 0 x1357 0 0.0207923249517024
Gyc1_1358 y1 0 x1358 0 -0.0314622224743914
Gyc1_1359 y1 0 x1359 0 0.0310802081089804
Gyc1_1360 y1 0 x1360 0 0.0216498808183829
Gyc1_1361 y1 0 x1361 0 -0.0937873388058954
Gyc1_1362 y1 0 x1362 0 0.079034802488912
Gyc1_1363 y1 0 x1363 0 -0.0266353754043708
Gyc1_1364 y1 0 x1364 0 0.0655981783982183
Gyc1_1365 y1 0 x1365 0 -0.0166341745995707
Gyc1_1366 y1 0 x1366 0 0.0128676819931694
Gyc1_1367 y1 0 x1367 0 0.00992631463445867
Gyc1_1368 y1 0 x1368 0 -0.046644477132823
Gyc1_1369 y1 0 x1369 0 -0.0145792957421774
Gyc1_1370 y1 0 x1370 0 -0.0196473274055042
Gyc1_1371 y1 0 x1371 0 0.0156689973739115
Gyc1_1372 y1 0 x1372 0 0.0291477049212213
Gyc1_1373 y1 0 x1373 0 -0.020361887508861
Gyc1_1374 y1 0 x1374 0 -0.0482893727887497
Gyc1_1375 y1 0 x1375 0 0.0167751888826163
Gyc1_1376 y1 0 x1376 0 0.041202955899886
Gyc1_1377 y1 0 x1377 0 0.0210255468834735
Gyc1_1378 y1 0 x1378 0 0.0296892678345895
Gyc1_1379 y1 0 x1379 0 -0.0347292420777175
Gyc1_1380 y1 0 x1380 0 -0.0374914123861875
Gyc1_1381 y1 0 x1381 0 0.0208242129288563
Gyc1_1382 y1 0 x1382 0 0.0374269616682147
Gyc1_1383 y1 0 x1383 0 0.00808764768740207
Gyc1_1384 y1 0 x1384 0 -0.024463660583131
Gyc1_1385 y1 0 x1385 0 -0.0168939158153349
Gyc1_1386 y1 0 x1386 0 -0.177204785429858
Gyc1_1387 y1 0 x1387 0 0.013962085470779
Gyc1_1388 y1 0 x1388 0 0.032649867990074
Gyc1_1389 y1 0 x1389 0 0.0248178423606218
Gyc1_1390 y1 0 x1390 0 -0.0216780065183514
Gyc1_1391 y1 0 x1391 0 -0.0252334550927795
Gyc1_1392 y1 0 x1392 0 0.0190941374440732
Gyc1_1393 y1 0 x1393 0 0.0272554399259301
Gyc1_1394 y1 0 x1394 0 0.0663355841388624
Gyc1_1395 y1 0 x1395 0 -0.0205302955402582
Gyc1_1396 y1 0 x1396 0 -0.0221772131008072
Gyc1_1397 y1 0 x1397 0 -0.0371077283165572
Gyc1_1398 y1 0 x1398 0 0.0306253349158099
Gyc1_1399 y1 0 x1399 0 -0.0312463601923977
Gyc1_1400 y1 0 x1400 0 0.0176127763905695
Gyc1_1401 y1 0 x1401 0 -0.0241984189524232
Gyc1_1402 y1 0 x1402 0 -0.0351871572145942
Gyc1_1403 y1 0 x1403 0 -0.00678397470770563
Gyc1_1404 y1 0 x1404 0 -0.028132466947539
Gyc1_1405 y1 0 x1405 0 0.0205011850622515
Gyc1_1406 y1 0 x1406 0 0.040838112757806
Gyc1_1407 y1 0 x1407 0 -0.0375079710978285
Gyc1_1408 y1 0 x1408 0 0.0257482677089626
Gyc1_1409 y1 0 x1409 0 -0.302962799761433
Gyc1_1410 y1 0 x1410 0 0.0138740301850867
Gyc1_1411 y1 0 x1411 0 -0.00396041781868457
Gyc1_1412 y1 0 x1412 0 0.0338808748136168
Gyc1_1413 y1 0 x1413 0 -0.0233972343753139
Gyc1_1414 y1 0 x1414 0 -0.0411555383223355
Gyc1_1415 y1 0 x1415 0 0.0466401592647162
Gyc1_1416 y1 0 x1416 0 -0.0313358826643722
Gyc1_1417 y1 0 x1417 0 -0.0197537809921147
Gyc1_1418 y1 0 x1418 0 -0.00844302817979178
Gyc1_1419 y1 0 x1419 0 0.0203556204456504
Gyc1_1420 y1 0 x1420 0 -0.0259887338008175
Gyc1_1421 y1 0 x1421 0 0.0284008227060007
Gyc1_1422 y1 0 x1422 0 -0.0310168506280793
Gyc1_1423 y1 0 x1423 0 0.0295390293183448
Gyc1_1424 y1 0 x1424 0 0.0432671105932941
Gyc1_1425 y1 0 x1425 0 -0.0952009222944763
Gyc1_1426 y1 0 x1426 0 -0.00552596536510028
Gyc1_1427 y1 0 x1427 0 -0.133797138700348
Gyc1_1428 y1 0 x1428 0 -0.0212072250558169
Gyc1_1429 y1 0 x1429 0 0.0524422447754649
Gyc1_1430 y1 0 x1430 0 0.0438532627327034
Gyc1_1431 y1 0 x1431 0 0.0459591747337298
Gyc1_1432 y1 0 x1432 0 0.0259089552629029
Gyc1_1433 y1 0 x1433 0 -0.00469824395624816
Gyc1_1434 y1 0 x1434 0 0.0644830662555481
Gyc1_1435 y1 0 x1435 0 0.0268079859846699
Gyc1_1436 y1 0 x1436 0 -0.0608340940020062
Gyc1_1437 y1 0 x1437 0 -0.0241921847995255
Gyc1_1438 y1 0 x1438 0 0.025233733830495
Gyc1_1439 y1 0 x1439 0 -0.0248502632326878
Gyc1_1440 y1 0 x1440 0 -0.0231836122888167
Gyc1_1441 y1 0 x1441 0 -0.0193486551498421
Gyc1_1442 y1 0 x1442 0 -0.0116282342758863
Gyc1_1443 y1 0 x1443 0 0.00854805099121288
Gyc1_1444 y1 0 x1444 0 -0.00517003983655636
Gyc1_1445 y1 0 x1445 0 0.0261471514693973
Gyc1_1446 y1 0 x1446 0 -0.0245307128285614
Gyc1_1447 y1 0 x1447 0 -0.0282576238438567
Gyc1_1448 y1 0 x1448 0 -0.0277150835601743
Gyc1_1449 y1 0 x1449 0 -0.0270362938607574
Gyc1_1450 y1 0 x1450 0 0.0327272315284753
Gyc1_1451 y1 0 x1451 0 -0.0254947030632868
Gyc1_1452 y1 0 x1452 0 -0.0205989518020538
Gyc1_1453 y1 0 x1453 0 -1
Gyc1_1454 y1 0 x1454 0 -0.0209463860364519
Gyc1_1455 y1 0 x1455 0 -0.0126461334811468
Gyc1_1456 y1 0 x1456 0 -0.0163133386887193
Gyc1_1457 y1 0 x1457 0 0.0330971449222107
Gyc1_1458 y1 0 x1458 0 -0.022603221252583
Gyc1_1459 y1 0 x1459 0 -0.0170597656698596
Gyc1_1460 y1 0 x1460 0 0.0136890946535958
Gyc1_1461 y1 0 x1461 0 0.260593758101848
Gyc1_1462 y1 0 x1462 0 -0.122498942067012
Gyc1_1463 y1 0 x1463 0 0.0226714488334525
Gyc1_1464 y1 0 x1464 0 0.0181148361018779
Gyc1_1465 y1 0 x1465 0 -0.00362232746181633
Gyc1_1466 y1 0 x1466 0 0.0161352051686175
Gyc1_1467 y1 0 x1467 0 -0.00356646407771472
Gyc1_1468 y1 0 x1468 0 -0.0220790858555284
Gyc1_1469 y1 0 x1469 0 0.0248809641519161
Gyc1_1470 y1 0 x1470 0 -0.0187243671474055
Gyc1_1471 y1 0 x1471 0 -0.0133624817969128
Gyc1_1472 y1 0 x1472 0 -0.0289352624943067
Gyc1_1473 y1 0 x1473 0 0.0302831872087606
Gyc1_1474 y1 0 x1474 0 -0.0214014749540041
Gyc1_1475 y1 0 x1475 0 -0.0260583605673438
Gyc1_1476 y1 0 x1476 0 0.0186739278176636
Gyc1_1477 y1 0 x1477 0 0.0242793319174556
Gyc1_1478 y1 0 x1478 0 0.0352975332349387
Gyc1_1479 y1 0 x1479 0 -0.0191264944158378
Gyc1_1480 y1 0 x1480 0 0.706575606243755
Gyc1_1481 y1 0 x1481 0 -0.0193361478607302
Gyc1_1482 y1 0 x1482 0 0.0221270102020579
Gyc1_1483 y1 0 x1483 0 -0.954291190816715
Gyc1_1484 y1 0 x1484 0 -0.0310204273447883
Gyc1_1485 y1 0 x1485 0 0.010037370115796
Gyc1_1486 y1 0 x1486 0 0.0101330613061208
Gyc1_1487 y1 0 x1487 0 0.0293683029811191
Gyc1_1488 y1 0 x1488 0 0.0303953539396224
Gyc1_1489 y1 0 x1489 0 -0.0656229081406126
Gyc1_1490 y1 0 x1490 0 0.0247074536987539
Gyc1_1491 y1 0 x1491 0 -0.0537611661241303
Gyc1_1492 y1 0 x1492 0 0.0273211624247025
Gyc1_1493 y1 0 x1493 0 -0.308577932355367
Gyc1_1494 y1 0 x1494 0 0.0255466315971921
Gyc1_1495 y1 0 x1495 0 0.0244525735880868
Gyc1_1496 y1 0 x1496 0 -0.0233076908075537
Gyc1_1497 y1 0 x1497 0 0.0892697325828824
Gyc1_1498 y1 0 x1498 0 0.00156328325565323
Gyc1_1499 y1 0 x1499 0 -0.0113287847723478
Gyc1_1500 y1 0 x1500 0 -0.0126292132986249
Gyc1_1501 y1 0 x1501 0 0.00224148663178152
Gyc1_1502 y1 0 x1502 0 0.0289479237683894
Gyc1_1503 y1 0 x1503 0 0.165781979219652
Gyc1_1504 y1 0 x1504 0 -0.0205018264876851
Gyc1_1505 y1 0 x1505 0 -0.0298768238030037
Gyc1_1506 y1 0 x1506 0 -0.0362793375745313
Gyc1_1507 y1 0 x1507 0 0.0342963529355439
Gyc1_1508 y1 0 x1508 0 -0.0373720220240639
Gyc1_1509 y1 0 x1509 0 0.0339979263871424
Gyc1_1510 y1 0 x1510 0 -0.0250455277658747
Gyc1_1511 y1 0 x1511 0 0.0505541288053004
Gyc1_1512 y1 0 x1512 0 0.653416059575291
Gyc1_1513 y1 0 x1513 0 -0.058528299683379
Gyc1_1514 y1 0 x1514 0 -0.0310149419960676
Gyc1_1515 y1 0 x1515 0 -0.00394498092162708
Gyc1_1516 y1 0 x1516 0 -0.0289672450923429
Gyc1_1517 y1 0 x1517 0 0.019459147470001
Gyc1_1518 y1 0 x1518 0 0.0128165769612177
Gyc1_1519 y1 0 x1519 0 -0.0264305919765579
Gyc1_1520 y1 0 x1520 0 -0.0199332396139606
Gyc1_1521 y1 0 x1521 0 0.0128559653257858
Gyc1_1522 y1 0 x1522 0 0.0785039884728083
Gyc1_1523 y1 0 x1523 0 0.0143020541034598
Gyc1_1524 y1 0 x1524 0 -0.00910374186958633
Gyc1_1525 y1 0 x1525 0 -0.00890840487352485
Gyc1_1526 y1 0 x1526 0 -0.0267139704617201
Gyc1_1527 y1 0 x1527 0 -0.034699016680192
Gyc1_1528 y1 0 x1528 0 0.00638932763054962
Gyc1_1529 y1 0 x1529 0 -0.00796240036596703
Gyc1_1530 y1 0 x1530 0 -0.0245189938952374
Gyc1_1531 y1 0 x1531 0 0.0287676856685556
Gyc1_1532 y1 0 x1532 0 -0.0313658626247588
Gyc1_1533 y1 0 x1533 0 0.0292956166317971
Gyc1_1534 y1 0 x1534 0 0.0331839965072001
Gyc1_1535 y1 0 x1535 0 0.0234924790858531
Gyc1_1536 y1 0 x1536 0 -0.0933749047828146
Gyc1_1537 y1 0 x1537 0 -0.00993297323695395
Gyc1_1538 y1 0 x1538 0 0.0199721611132404
Gyc1_1539 y1 0 x1539 0 0.0202147123453211
Gyc1_1540 y1 0 x1540 0 0.0343758410501239
Gyc1_1541 y1 0 x1541 0 0.0337222252967354
Gyc1_1542 y1 0 x1542 0 -0.0110940435217057
Gyc1_1543 y1 0 x1543 0 -0.0265671643756131
Gyc1_1544 y1 0 x1544 0 -0.0217766979378518
Gyc1_1545 y1 0 x1545 0 0.0111077748817256
Gyc1_1546 y1 0 x1546 0 -0.0287559784578905
Gyc1_1547 y1 0 x1547 0 -0.0233002720552533
Gyc1_1548 y1 0 x1548 0 -0.0293265769772924
Gyc1_1549 y1 0 x1549 0 0.0196867980234338
Gyc1_1550 y1 0 x1550 0 -0.0258161189330652
Gyc1_1551 y1 0 x1551 0 1
Gyc1_1552 y1 0 x1552 0 -0.026373028154591
Gyc1_1553 y1 0 x1553 0 -0.0210558412590185
Gyc1_1554 y1 0 x1554 0 -0.0172812524854833
Gyc1_1555 y1 0 x1555 0 0.0617760128261759
Gyc1_1556 y1 0 x1556 0 0.0262441749135716
Gyc1_1557 y1 0 x1557 0 -0.0135382306693118
Gyc1_1558 y1 0 x1558 0 0.0390193903519931
Gyc1_1559 y1 0 x1559 0 0.0220907210697965
Gyc1_1560 y1 0 x1560 0 0.0190594894891981
Gyc1_1561 y1 0 x1561 0 -0.0634218055118851
Gyc1_1562 y1 0 x1562 0 0.00405633233285839
Gyc1_1563 y1 0 x1563 0 -0.0109619148856904
Gyc1_1564 y1 0 x1564 0 -0.0319168334045588
Gyc1_1565 y1 0 x1565 0 -0.0346050218165637
Gyc1_1566 y1 0 x1566 0 0.0130832318653254
Gyc1_1567 y1 0 x1567 0 0.0281813637881807
Gyc1_1568 y1 0 x1568 0 -0.0564811689213441
Gyc1_1569 y1 0 x1569 0 0.0223733383339309
Gyc1_1570 y1 0 x1570 0 0.0204808537988391
Gyc1_1571 y1 0 x1571 0 -0.0268671178040414
Gyc1_1572 y1 0 x1572 0 0.0334586521271445
Gyc1_1573 y1 0 x1573 0 0.0229714587005257
Gyc1_1574 y1 0 x1574 0 0.0334785498995261
Gyc1_1575 y1 0 x1575 0 0.0407968888068999
Gyc1_1576 y1 0 x1576 0 0.1142158769969
Gyc1_1577 y1 0 x1577 0 0.0352322181897299
Gyc1_1578 y1 0 x1578 0 -0.0127740700345019
Gyc1_1579 y1 0 x1579 0 0.0139804880693943
Gyc1_1580 y1 0 x1580 0 0.0396526475912192
Gyc1_1581 y1 0 x1581 0 0.0421423111476503
Gyc1_1582 y1 0 x1582 0 0.0250208451112281
Gyc1_1583 y1 0 x1583 0 0.0311846921520738
Gyc1_1584 y1 0 x1584 0 0.0184119083993307
Gyc1_1585 y1 0 x1585 0 -0.00205764962253491
Gyc1_1586 y1 0 x1586 0 0.0272931987348298
Gyc1_1587 y1 0 x1587 0 -0.0420804368998569
Gyc1_1588 y1 0 x1588 0 0.0173298161170755
Gyc1_1589 y1 0 x1589 0 -0.0251793511894766
Gyc1_1590 y1 0 x1590 0 -0.0249580686053487
Gyc1_1591 y1 0 x1591 0 0.0762261509270341
Gyc1_1592 y1 0 x1592 0 -0.0200816538153769
Gyc1_1593 y1 0 x1593 0 -0.0405655270730253
Gyc1_1594 y1 0 x1594 0 0.0368231521982465
Gyc1_1595 y1 0 x1595 0 0.0405997677089457
Gyc1_1596 y1 0 x1596 0 -0.0269979791853058
Gyc1_1597 y1 0 x1597 0 -0.0246380331594294
Gyc1_1598 y1 0 x1598 0 0.00681919079905246
Gyc1_1599 y1 0 x1599 0 0.0074706424937459
Gyc1_1600 y1 0 x1600 0 0.0138461318865105
Gyc1_1601 y1 0 x1601 0 0.0248459856969482
Gyc1_1602 y1 0 x1602 0 -0.335467963528222
Gyc2_1 y2 0 x1 0 -0.0613095722658684
Gyc2_2 y2 0 x2 0 0.0608593408467446
Gyc2_3 y2 0 x3 0 -0.0499680517101837
Gyc2_4 y2 0 x4 0 -0.0820447482219613
Gyc2_5 y2 0 x5 0 -0.0617652199166415
Gyc2_6 y2 0 x6 0 0.165728517107174
Gyc2_7 y2 0 x7 0 0.159378880082134
Gyc2_8 y2 0 x8 0 -0.044147105007466
Gyc2_9 y2 0 x9 0 0.0954927124366981
Gyc2_10 y2 0 x10 0 0.117400515290567
Gyc2_11 y2 0 x11 0 0.15628181026714
Gyc2_12 y2 0 x12 0 0.0861757853343058
Gyc2_13 y2 0 x13 0 -0.218308920693104
Gyc2_14 y2 0 x14 0 0.0656666008826586
Gyc2_15 y2 0 x15 0 -0.0236226351550356
Gyc2_16 y2 0 x16 0 0.0974366470745647
Gyc2_17 y2 0 x17 0 -0.0696929191632578
Gyc2_18 y2 0 x18 0 -0.361636404594711
Gyc2_19 y2 0 x19 0 0.0520204880473498
Gyc2_20 y2 0 x20 0 0.118136019735881
Gyc2_21 y2 0 x21 0 -0.0282094420564341
Gyc2_22 y2 0 x22 0 -0.155506184240109
Gyc2_23 y2 0 x23 0 -0.0944570341632054
Gyc2_24 y2 0 x24 0 -0.113107435927873
Gyc2_25 y2 0 x25 0 -0.138424176771755
Gyc2_26 y2 0 x26 0 0.0556847732869524
Gyc2_27 y2 0 x27 0 -0.51697517329734
Gyc2_28 y2 0 x28 0 0.0747804020134338
Gyc2_29 y2 0 x29 0 -0.129913453308786
Gyc2_30 y2 0 x30 0 0.0514154564706046
Gyc2_31 y2 0 x31 0 -0.123792945941594
Gyc2_32 y2 0 x32 0 0.0480405412172027
Gyc2_33 y2 0 x33 0 -0.0955100153911476
Gyc2_34 y2 0 x34 0 -0.0208455203135179
Gyc2_35 y2 0 x35 0 0.01902434334897
Gyc2_36 y2 0 x36 0 -0.0999123520600306
Gyc2_37 y2 0 x37 0 0.0987699115672825
Gyc2_38 y2 0 x38 0 -0.0257324685895143
Gyc2_39 y2 0 x39 0 0.0841154594807846
Gyc2_40 y2 0 x40 0 1
Gyc2_41 y2 0 x41 0 -0.149314062342692
Gyc2_42 y2 0 x42 0 0.0580921859662313
Gyc2_43 y2 0 x43 0 -0.0842020907185935
Gyc2_44 y2 0 x44 0 0.102209318235911
Gyc2_45 y2 0 x45 0 -0.0940982623692445
Gyc2_46 y2 0 x46 0 -0.0980900040333489
Gyc2_47 y2 0 x47 0 -0.0510090422939495
Gyc2_48 y2 0 x48 0 -0.189029707089411
Gyc2_49 y2 0 x49 0 -0.416972305955835
Gyc2_50 y2 0 x50 0 0.112256234550292
Gyc2_51 y2 0 x51 0 0.0263350621023178
Gyc2_52 y2 0 x52 0 0.126811021394714
Gyc2_53 y2 0 x53 0 -0.159103694279122
Gyc2_54 y2 0 x54 0 0.0901201693413958
Gyc2_55 y2 0 x55 0 -0.0922062902197064
Gyc2_56 y2 0 x56 0 -0.0411313102371984
Gyc2_57 y2 0 x57 0 0.105432843586274
Gyc2_58 y2 0 x58 0 -0.031507715779932
Gyc2_59 y2 0 x59 0 -0.0450926174310101
Gyc2_60 y2 0 x60 0 -0.113655692013565
Gyc2_61 y2 0 x61 0 1
Gyc2_62 y2 0 x62 0 -0.13550276141074
Gyc2_63 y2 0 x63 0 -0.00686438931446288
Gyc2_64 y2 0 x64 0 0.0763140962740398
Gyc2_65 y2 0 x65 0 0.000707338079352287
Gyc2_66 y2 0 x66 0 0.0864340447247554
Gyc2_67 y2 0 x67 0 -0.127631813224265
Gyc2_68 y2 0 x68 0 -0.02988045279323
Gyc2_69 y2 0 x69 0 -0.0660713253630543
Gyc2_70 y2 0 x70 0 -0.159349180624713
Gyc2_71 y2 0 x71 0 -0.0252008901910511
Gyc2_72 y2 0 x72 0 -0.12884023544172
Gyc2_73 y2 0 x73 0 0.116873044114598
Gyc2_74 y2 0 x74 0 -0.115077646029385
Gyc2_75 y2 0 x75 0 -0.0161296333448569
Gyc2_76 y2 0 x76 0 -0.102804863541921
Gyc2_77 y2 0 x77 0 0.0807836595226542
Gyc2_78 y2 0 x78 0 0.169987540413966
Gyc2_79 y2 0 x79 0 -0.313811043562439
Gyc2_80 y2 0 x80 0 0.082338026869269
Gyc2_81 y2 0 x81 0 -0.0780836438999335
Gyc2_82 y2 0 x82 0 -0.18500220660266
Gyc2_83 y2 0 x83 0 -0.0485612775394968
Gyc2_84 y2 0 x84 0 -0.24078118614963
Gyc2_85 y2 0 x85 0 0.0404721417762776
Gyc2_86 y2 0 x86 0 0.0830000070959385
Gyc2_87 y2 0 x87 0 0.567414585446288
Gyc2_88 y2 0 x88 0 -0.0991195572270392
Gyc2_89 y2 0 x89 0 0.108619740906346
Gyc2_90 y2 0 x90 0 0.423213092144238
Gyc2_91 y2 0 x91 0 0.0823166399682088
Gyc2_92 y2 0 x92 0 1
Gyc2_93 y2 0 x93 0 0.153497297578711
Gyc2_94 y2 0 x94 0 -0.0620457381107954
Gyc2_95 y2 0 x95 0 -0.0866234719342059
Gyc2_96 y2 0 x96 0 -0.239202118252329
Gyc2_97 y2 0 x97 0 -0.0267973071687741
Gyc2_98 y2 0 x98 0 -0.101511476562871
Gyc2_99 y2 0 x99 0 -0.0666645837182702
Gyc2_100 y2 0 x100 0 -0.25471954034551
Gyc2_101 y2 0 x101 0 -0.0474372384549574
Gyc2_102 y2 0 x102 0 -0.129704347221314
Gyc2_103 y2 0 x103 0 0.00315207877350674
Gyc2_104 y2 0 x104 0 -0.10797009985105
Gyc2_105 y2 0 x105 0 0.112809659893888
Gyc2_106 y2 0 x106 0 -0.0288074386441916
Gyc2_107 y2 0 x107 0 0.104128334184867
Gyc2_108 y2 0 x108 0 -0.00501270700871351
Gyc2_109 y2 0 x109 0 -0.0237044495750154
Gyc2_110 y2 0 x110 0 -0.10734581489883
Gyc2_111 y2 0 x111 0 0.108020041184784
Gyc2_112 y2 0 x112 0 -0.0913953370153456
Gyc2_113 y2 0 x113 0 0.175075457944276
Gyc2_114 y2 0 x114 0 -0.0923865149863592
Gyc2_115 y2 0 x115 0 0.0841097315054589
Gyc2_116 y2 0 x116 0 0.22443269728167
Gyc2_117 y2 0 x117 0 0.0574004194233827
Gyc2_118 y2 0 x118 0 0.131834986008329
Gyc2_119 y2 0 x119 0 0.0908838156267204
Gyc2_120 y2 0 x120 0 0.130874090266709
Gyc2_121 y2 0 x121 0 -0.0599852119566297
Gyc2_122 y2 0 x122 0 -0.128397211709396
Gyc2_123 y2 0 x123 0 -0.205415453104912
Gyc2_124 y2 0 x124 0 0.0709475337495983
Gyc2_125 y2 0 x125 0 -0.0511492494222286
Gyc2_126 y2 0 x126 0 -0.12783554736382
Gyc2_127 y2 0 x127 0 -0.0419664095056249
Gyc2_128 y2 0 x128 0 -0.122212708605017
Gyc2_129 y2 0 x129 0 -0.113012579691365
Gyc2_130 y2 0 x130 0 0.0255379848456497
Gyc2_131 y2 0 x131 0 -0.135662551042328
Gyc2_132 y2 0 x132 0 0.104571957854092
Gyc2_133 y2 0 x133 0 0.101488173526922
Gyc2_134 y2 0 x134 0 -0.0536298396292153
Gyc2_135 y2 0 x135 0 -0.0847467974841788
Gyc2_136 y2 0 x136 0 -0.161412671761843
Gyc2_137 y2 0 x137 0 0.103505669185963
Gyc2_138 y2 0 x138 0 -0.0721518770019033
Gyc2_139 y2 0 x139 0 0.123127617022541
Gyc2_140 y2 0 x140 0 0.0725310227508353
Gyc2_141 y2 0 x141 0 -0.0457289044486992
Gyc2_142 y2 0 x142 0 -0.112541212377217
Gyc2_143 y2 0 x143 0 -0.115401479772214
Gyc2_144 y2 0 x144 0 0.0574137223439544
Gyc2_145 y2 0 x145 0 0.0787505262111815
Gyc2_146 y2 0 x146 0 0.227175247624844
Gyc2_147 y2 0 x147 0 1
Gyc2_148 y2 0 x148 0 -0.101718986432168
Gyc2_149 y2 0 x149 0 -0.0771520464215817
Gyc2_150 y2 0 x150 0 -0.291637450620385
Gyc2_151 y2 0 x151 0 -0.101008080833122
Gyc2_152 y2 0 x152 0 0.0304247154156433
Gyc2_153 y2 0 x153 0 -0.0948370065511739
Gyc2_154 y2 0 x154 0 0.0286909167373701
Gyc2_155 y2 0 x155 0 0.0664169214532511
Gyc2_156 y2 0 x156 0 0.13207300971824
Gyc2_157 y2 0 x157 0 0.849621783352601
Gyc2_158 y2 0 x158 0 -0.0720862748093391
Gyc2_159 y2 0 x159 0 0.618081710472809
Gyc2_160 y2 0 x160 0 -1
Gyc2_161 y2 0 x161 0 -0.199416430334962
Gyc2_162 y2 0 x162 0 0.0770170865945222
Gyc2_163 y2 0 x163 0 -0.0726623214714648
Gyc2_164 y2 0 x164 0 -0.116475906727983
Gyc2_165 y2 0 x165 0 -0.00832585301165825
Gyc2_166 y2 0 x166 0 -0.205450199915595
Gyc2_167 y2 0 x167 0 -0.153218332261428
Gyc2_168 y2 0 x168 0 0.0927428170120762
Gyc2_169 y2 0 x169 0 0.102133883114662
Gyc2_170 y2 0 x170 0 -0.0916196400640586
Gyc2_171 y2 0 x171 0 0.0599385497820557
Gyc2_172 y2 0 x172 0 0.153098418074561
Gyc2_173 y2 0 x173 0 -0.0882578758424172
Gyc2_174 y2 0 x174 0 -0.121140463130983
Gyc2_175 y2 0 x175 0 0.0784722869716771
Gyc2_176 y2 0 x176 0 0.120067584023267
Gyc2_177 y2 0 x177 0 -0.129572559755673
Gyc2_178 y2 0 x178 0 0.0771132105861104
Gyc2_179 y2 0 x179 0 0.102067087619253
Gyc2_180 y2 0 x180 0 -0.0762711560804404
Gyc2_181 y2 0 x181 0 -0.197631209119129
Gyc2_182 y2 0 x182 0 -0.781394957833461
Gyc2_183 y2 0 x183 0 0.11749931544045
Gyc2_184 y2 0 x184 0 -0.130027615349558
Gyc2_185 y2 0 x185 0 0.114883876170668
Gyc2_186 y2 0 x186 0 -0.0904729593659939
Gyc2_187 y2 0 x187 0 -0.0850231319911251
Gyc2_188 y2 0 x188 0 -0.187414265721487
Gyc2_189 y2 0 x189 0 -0.0865530379525283
Gyc2_190 y2 0 x190 0 -0.175141172039246
Gyc2_191 y2 0 x191 0 -0.0310832248592483
Gyc2_192 y2 0 x192 0 -0.0957078358053966
Gyc2_193 y2 0 x193 0 0.0753435995556787
Gyc2_194 y2 0 x194 0 0.118375036757282
Gyc2_195 y2 0 x195 0 0.209848361931312
Gyc2_196 y2 0 x196 0 -0.0958665509045329
Gyc2_197 y2 0 x197 0 -0.0855329868307132
Gyc2_198 y2 0 x198 0 -0.0213898550261229
Gyc2_199 y2 0 x199 0 -0.0864320109496864
Gyc2_200 y2 0 x200 0 -0.220871727013267
Gyc2_201 y2 0 x201 0 0.193744031909729
Gyc2_202 y2 0 x202 0 0.10105969220689
Gyc2_203 y2 0 x203 0 -0.0981042645307734
Gyc2_204 y2 0 x204 0 0.0452781724145052
Gyc2_205 y2 0 x205 0 -0.462466198927902
Gyc2_206 y2 0 x206 0 -0.000382466200414262
Gyc2_207 y2 0 x207 0 0.11764917792258
Gyc2_208 y2 0 x208 0 -0.577920013242202
Gyc2_209 y2 0 x209 0 -0.0583268416820292
Gyc2_210 y2 0 x210 0 -0.0957604163190847
Gyc2_211 y2 0 x211 0 -1
Gyc2_212 y2 0 x212 0 0.815554137088267
Gyc2_213 y2 0 x213 0 -0.102064446136013
Gyc2_214 y2 0 x214 0 -0.0830313319305245
Gyc2_215 y2 0 x215 0 -0.0951128602475109
Gyc2_216 y2 0 x216 0 0.0590729626452356
Gyc2_217 y2 0 x217 0 -0.0715960593632247
Gyc2_218 y2 0 x218 0 -0.0952999063972793
Gyc2_219 y2 0 x219 0 -0.110769078424412
Gyc2_220 y2 0 x220 0 0.0679987203523252
Gyc2_221 y2 0 x221 0 0.191868765510806
Gyc2_222 y2 0 x222 0 -0.0678095077157542
Gyc2_223 y2 0 x223 0 0.105177415137935
Gyc2_224 y2 0 x224 0 -0.0811881577246942
Gyc2_225 y2 0 x225 0 0.308435415760536
Gyc2_226 y2 0 x226 0 0.290530022281069
Gyc2_227 y2 0 x227 0 0.078904755420201
Gyc2_228 y2 0 x228 0 -0.0486097425494303
Gyc2_229 y2 0 x229 0 0.106602171426817
Gyc2_230 y2 0 x230 0 -0.124812823983669
Gyc2_231 y2 0 x231 0 -0.0740907286395171
Gyc2_232 y2 0 x232 0 0.117023970718932
Gyc2_233 y2 0 x233 0 0.012114530202548
Gyc2_234 y2 0 x234 0 0.0551023327473222
Gyc2_235 y2 0 x235 0 -0.0548440021254164
Gyc2_236 y2 0 x236 0 -0.875169060778351
Gyc2_237 y2 0 x237 0 -0.097613534387124
Gyc2_238 y2 0 x238 0 0.0397939261504303
Gyc2_239 y2 0 x239 0 -0.114362793522258
Gyc2_240 y2 0 x240 0 -0.128364631859552
Gyc2_241 y2 0 x241 0 -0.121930962082854
Gyc2_242 y2 0 x242 0 0.0774848203234099
Gyc2_243 y2 0 x243 0 -0.119191257243948
Gyc2_244 y2 0 x244 0 0.201086737886786
Gyc2_245 y2 0 x245 0 0.800163754621766
Gyc2_246 y2 0 x246 0 -0.0544475408637474
Gyc2_247 y2 0 x247 0 0.174025987299421
Gyc2_248 y2 0 x248 0 0.0886490659999472
Gyc2_249 y2 0 x249 0 -0.0673708521167617
Gyc2_250 y2 0 x250 0 -0.0957681608768778
Gyc2_251 y2 0 x251 0 0.556102706401893
Gyc2_252 y2 0 x252 0 0.0907444351382341
Gyc2_253 y2 0 x253 0 -0.0471711079370357
Gyc2_254 y2 0 x254 0 0.171535735822387
Gyc2_255 y2 0 x255 0 0.122946823176413
Gyc2_256 y2 0 x256 0 -0.100322416836891
Gyc2_257 y2 0 x257 0 -0.104356616160329
Gyc2_258 y2 0 x258 0 -0.0994884547231786
Gyc2_259 y2 0 x259 0 0.058645855481652
Gyc2_260 y2 0 x260 0 -0.0994805339550955
Gyc2_261 y2 0 x261 0 0.0774666988915637
Gyc2_262 y2 0 x262 0 -0.206509524520517
Gyc2_263 y2 0 x263 0 -0.0354346468036905
Gyc2_264 y2 0 x264 0 -0.0754632317592863
Gyc2_265 y2 0 x265 0 -0.0607943280280388
Gyc2_266 y2 0 x266 0 0.0461689056480666
Gyc2_267 y2 0 x267 0 -0.00595624701121563
Gyc2_268 y2 0 x268 0 0.0520352483764552
Gyc2_269 y2 0 x269 0 0.121461874419156
Gyc2_270 y2 0 x270 0 0.0483650808606929
Gyc2_271 y2 0 x271 0 0.034245692972357
Gyc2_272 y2 0 x272 0 0.0102530227719455
Gyc2_273 y2 0 x273 0 -0.00785975683343191
Gyc2_274 y2 0 x274 0 0.0563032537899998
Gyc2_275 y2 0 x275 0 -0.0509398806947516
Gyc2_276 y2 0 x276 0 -0.0373957747624223
Gyc2_277 y2 0 x277 0 0.010629897433525
Gyc2_278 y2 0 x278 0 -0.0856575561543449
Gyc2_279 y2 0 x279 0 0.141293636212033
Gyc2_280 y2 0 x280 0 0.00134991356510416
Gyc2_281 y2 0 x281 0 0.0876082010326971
Gyc2_282 y2 0 x282 0 -0.0636228092712534
Gyc2_283 y2 0 x283 0 0.0488985821811735
Gyc2_284 y2 0 x284 0 -0.00203585130001215
Gyc2_285 y2 0 x285 0 0.0973639068097899
Gyc2_286 y2 0 x286 0 -0.0505019252276504
Gyc2_287 y2 0 x287 0 -0.0763984317726781
Gyc2_288 y2 0 x288 0 0.304973018120646
Gyc2_289 y2 0 x289 0 -0.0395636470626578
Gyc2_290 y2 0 x290 0 0.0183570319022618
Gyc2_291 y2 0 x291 0 0.0717660848303957
Gyc2_292 y2 0 x292 0 0.125955096335396
Gyc2_293 y2 0 x293 0 0.0334643960747404
Gyc2_294 y2 0 x294 0 -0.0537347004064339
Gyc2_295 y2 0 x295 0 -0.0429662596319135
Gyc2_296 y2 0 x296 0 0.0521964787682661
Gyc2_297 y2 0 x297 0 -0.173824255020819
Gyc2_298 y2 0 x298 0 0.108608081073527
Gyc2_299 y2 0 x299 0 -0.0310327387512892
Gyc2_300 y2 0 x300 0 -0.163124570944896
Gyc2_301 y2 0 x301 0 -0.00950765850281034
Gyc2_302 y2 0 x302 0 -0.0446181100466772
Gyc2_303 y2 0 x303 0 0.0704896854557916
Gyc2_304 y2 0 x304 0 0.153815915423508
Gyc2_305 y2 0 x305 0 0.0646199045804458
Gyc2_306 y2 0 x306 0 0.132875613439886
Gyc2_307 y2 0 x307 0 0.0964465021201247
Gyc2_308 y2 0 x308 0 0.0177477039329335
Gyc2_309 y2 0 x309 0 -0.0722213317149636
Gyc2_310 y2 0 x310 0 -0.134630862950794
Gyc2_311 y2 0 x311 0 -0.0600432252293942
Gyc2_312 y2 0 x312 0 0.0802387105792
Gyc2_313 y2 0 x313 0 -1
Gyc2_314 y2 0 x314 0 0.0846717211909411
Gyc2_315 y2 0 x315 0 0.0298321084511859
Gyc2_316 y2 0 x316 0 0.0863706623239656
Gyc2_317 y2 0 x317 0 -0.109405574174544
Gyc2_318 y2 0 x318 0 -0.170446612967699
Gyc2_319 y2 0 x319 0 -0.407589312497056
Gyc2_320 y2 0 x320 0 0.0919527077274289
Gyc2_321 y2 0 x321 0 0.0539722408645452
Gyc2_322 y2 0 x322 0 0.113638387397771
Gyc2_323 y2 0 x323 0 0.00789537247808374
Gyc2_324 y2 0 x324 0 -0.0505764467373434
Gyc2_325 y2 0 x325 0 -0.0589623972375951
Gyc2_326 y2 0 x326 0 0.0649520622792522
Gyc2_327 y2 0 x327 0 0.0515258601807503
Gyc2_328 y2 0 x328 0 0.109169653585962
Gyc2_329 y2 0 x329 0 0.0439739637070596
Gyc2_330 y2 0 x330 0 0.0898877371509969
Gyc2_331 y2 0 x331 0 0.113691468809004
Gyc2_332 y2 0 x332 0 0.434373307085526
Gyc2_333 y2 0 x333 0 -0.0141615097738694
Gyc2_334 y2 0 x334 0 0.21048955378403
Gyc2_335 y2 0 x335 0 0.0207368729639311
Gyc2_336 y2 0 x336 0 0.119049921559307
Gyc2_337 y2 0 x337 0 -0.040965049810528
Gyc2_338 y2 0 x338 0 -0.0445336494978117
Gyc2_339 y2 0 x339 0 -0.0114879910622027
Gyc2_340 y2 0 x340 0 -0.110471847020386
Gyc2_341 y2 0 x341 0 -0.0188706256408354
Gyc2_342 y2 0 x342 0 -0.107161176913876
Gyc2_343 y2 0 x343 0 0.0867239714904413
Gyc2_344 y2 0 x344 0 0.0973987865866658
Gyc2_345 y2 0 x345 0 0.059592386761632
Gyc2_346 y2 0 x346 0 0.121292764744656
Gyc2_347 y2 0 x347 0 -0.199203494566676
Gyc2_348 y2 0 x348 0 0.0617527237238577
Gyc2_349 y2 0 x349 0 0.0639523457415923
Gyc2_350 y2 0 x350 0 0.120955253825155
Gyc2_351 y2 0 x351 0 -0.066396822606291
Gyc2_352 y2 0 x352 0 -0.0082514510616765
Gyc2_353 y2 0 x353 0 0.0734723856564427
Gyc2_354 y2 0 x354 0 0.451376995634544
Gyc2_355 y2 0 x355 0 -0.00411606833605489
Gyc2_356 y2 0 x356 0 -0.109043601167611
Gyc2_357 y2 0 x357 0 0.0693601094627055
Gyc2_358 y2 0 x358 0 -0.103620020727423
Gyc2_359 y2 0 x359 0 -0.0636556092299659
Gyc2_360 y2 0 x360 0 0.118466477290491
Gyc2_361 y2 0 x361 0 -1
Gyc2_362 y2 0 x362 0 -0.190868326822189
Gyc2_363 y2 0 x363 0 -0.131460392422118
Gyc2_364 y2 0 x364 0 0.100905599746807
Gyc2_365 y2 0 x365 0 0.0591342786368174
Gyc2_366 y2 0 x366 0 0.106178230707311
Gyc2_367 y2 0 x367 0 -0.106737115824822
Gyc2_368 y2 0 x368 0 -0.118245463377419
Gyc2_369 y2 0 x369 0 -0.102167200239761
Gyc2_370 y2 0 x370 0 -0.124713072454316
Gyc2_371 y2 0 x371 0 0.0828539624920359
Gyc2_372 y2 0 x372 0 0.140266884726928
Gyc2_373 y2 0 x373 0 0.104829246666843
Gyc2_374 y2 0 x374 0 1
Gyc2_375 y2 0 x375 0 0.0941992500720495
Gyc2_376 y2 0 x376 0 0.0346297822989133
Gyc2_377 y2 0 x377 0 -0.138002764078367
Gyc2_378 y2 0 x378 0 0.0877931852797204
Gyc2_379 y2 0 x379 0 -0.104571588246142
Gyc2_380 y2 0 x380 0 -0.190723851106781
Gyc2_381 y2 0 x381 0 0.625035365964299
Gyc2_382 y2 0 x382 0 0.123198690560271
Gyc2_383 y2 0 x383 0 0.121791334823007
Gyc2_384 y2 0 x384 0 -0.0933291026765511
Gyc2_385 y2 0 x385 0 -0.100153558980193
Gyc2_386 y2 0 x386 0 0.104854224536547
Gyc2_387 y2 0 x387 0 -0.101227473847795
Gyc2_388 y2 0 x388 0 0.0302121136121176
Gyc2_389 y2 0 x389 0 -0.153487944647354
Gyc2_390 y2 0 x390 0 -0.104042636298881
Gyc2_391 y2 0 x391 0 0.0870068455398906
Gyc2_392 y2 0 x392 0 -0.09118680238975
Gyc2_393 y2 0 x393 0 -0.104264132220686
Gyc2_394 y2 0 x394 0 -0.11215081047685
Gyc2_395 y2 0 x395 0 0.0316769251546212
Gyc2_396 y2 0 x396 0 0.102039097873326
Gyc2_397 y2 0 x397 0 -0.0864944101074042
Gyc2_398 y2 0 x398 0 -0.116180621549808
Gyc2_399 y2 0 x399 0 -0.0913681980248923
Gyc2_400 y2 0 x400 0 0.114669011111972
Gyc2_401 y2 0 x401 0 0.12610999069163
Gyc2_402 y2 0 x402 0 -0.0560380884680846
Gyc2_403 y2 0 x403 0 0.118929008275636
Gyc2_404 y2 0 x404 0 -0.0472888416638188
Gyc2_405 y2 0 x405 0 0.0936710868283271
Gyc2_406 y2 0 x406 0 0.0762486150612961
Gyc2_407 y2 0 x407 0 -0.141056154503961
Gyc2_408 y2 0 x408 0 0.116536273015726
Gyc2_409 y2 0 x409 0 0.0824105449686586
Gyc2_410 y2 0 x410 0 0.0102123685162933
Gyc2_411 y2 0 x411 0 0.298029439251091
Gyc2_412 y2 0 x412 0 0.105726269438233
Gyc2_413 y2 0 x413 0 0.0820359503035985
Gyc2_414 y2 0 x414 0 -0.233950770445262
Gyc2_415 y2 0 x415 0 0.0851615946780369
Gyc2_416 y2 0 x416 0 0.102186953016143
Gyc2_417 y2 0 x417 0 -0.107518688851899
Gyc2_418 y2 0 x418 0 -0.061877680612676
Gyc2_419 y2 0 x419 0 -0.585644482144753
Gyc2_420 y2 0 x420 0 -0.128875966805034
Gyc2_421 y2 0 x421 0 0.0490255768836665
Gyc2_422 y2 0 x422 0 -0.21692216985828
Gyc2_423 y2 0 x423 0 -1
Gyc2_424 y2 0 x424 0 -0.160993117734202
Gyc2_425 y2 0 x425 0 0.0725854294109366
Gyc2_426 y2 0 x426 0 -0.0818872552338405
Gyc2_427 y2 0 x427 0 0.0701415662657309
Gyc2_428 y2 0 x428 0 -0.0853701391414569
Gyc2_429 y2 0 x429 0 0.116182635343798
Gyc2_430 y2 0 x430 0 -0.0832149694234709
Gyc2_431 y2 0 x431 0 -0.0692970154229934
Gyc2_432 y2 0 x432 0 -0.0947867745177131
Gyc2_433 y2 0 x433 0 0.0803678426768832
Gyc2_434 y2 0 x434 0 -0.0594539384736751
Gyc2_435 y2 0 x435 0 0.078480583653126
Gyc2_436 y2 0 x436 0 -0.0151492078764308
Gyc2_437 y2 0 x437 0 -0.0605263793240284
Gyc2_438 y2 0 x438 0 0.0771977317482436
Gyc2_439 y2 0 x439 0 0.0673186624444672
Gyc2_440 y2 0 x440 0 -0.0542487368287181
Gyc2_441 y2 0 x441 0 0.0659439818642684
Gyc2_442 y2 0 x442 0 0.0795572349920784
Gyc2_443 y2 0 x443 0 -0.0594234574461591
Gyc2_444 y2 0 x444 0 -0.0845966319705547
Gyc2_445 y2 0 x445 0 -0.0177099817522075
Gyc2_446 y2 0 x446 0 -0.0717901168954467
Gyc2_447 y2 0 x447 0 0.0912067905729694
Gyc2_448 y2 0 x448 0 0.0863587624568299
Gyc2_449 y2 0 x449 0 -0.105605790740065
Gyc2_450 y2 0 x450 0 0.0842233707349403
Gyc2_451 y2 0 x451 0 -0.028406281219011
Gyc2_452 y2 0 x452 0 0.0690410693498696
Gyc2_453 y2 0 x453 0 -0.13110429598298
Gyc2_454 y2 0 x454 0 0.0830802690471685
Gyc2_455 y2 0 x455 0 -0.0912393237300258
Gyc2_456 y2 0 x456 0 -0.853552325233326
Gyc2_457 y2 0 x457 0 0.286137095655868
Gyc2_458 y2 0 x458 0 -0.0863478426831149
Gyc2_459 y2 0 x459 0 -0.0976466719793945
Gyc2_460 y2 0 x460 0 -0.121099999369762
Gyc2_461 y2 0 x461 0 0.22101327910424
Gyc2_462 y2 0 x462 0 -0.00551496268536382
Gyc2_463 y2 0 x463 0 0.0429337940016587
Gyc2_464 y2 0 x464 0 0.18551195673412
Gyc2_465 y2 0 x465 0 0.0346629237564074
Gyc2_466 y2 0 x466 0 -0.0556548560744373
Gyc2_467 y2 0 x467 0 0.00843397130907148
Gyc2_468 y2 0 x468 0 0.0754311499552499
Gyc2_469 y2 0 x469 0 -0.135246388946615
Gyc2_470 y2 0 x470 0 0.0577778220104356
Gyc2_471 y2 0 x471 0 -0.0232275016903013
Gyc2_472 y2 0 x472 0 -0.0862524452946439
Gyc2_473 y2 0 x473 0 0.149669251192231
Gyc2_474 y2 0 x474 0 -0.0814638807545107
Gyc2_475 y2 0 x475 0 0.0739416289554796
Gyc2_476 y2 0 x476 0 -0.0369656710582866
Gyc2_477 y2 0 x477 0 0.141533328942614
Gyc2_478 y2 0 x478 0 -0.0654748510278281
Gyc2_479 y2 0 x479 0 0.0261142374232141
Gyc2_480 y2 0 x480 0 -0.0792933599655197
Gyc2_481 y2 0 x481 0 0.609723175591403
Gyc2_482 y2 0 x482 0 -0.10992877000533
Gyc2_483 y2 0 x483 0 0.0921682684916572
Gyc2_484 y2 0 x484 0 0.153072804971136
Gyc2_485 y2 0 x485 0 -0.191092062789632
Gyc2_486 y2 0 x486 0 -0.64833739845829
Gyc2_487 y2 0 x487 0 -0.128873219011012
Gyc2_488 y2 0 x488 0 -0.106037188350463
Gyc2_489 y2 0 x489 0 0.111935292371884
Gyc2_490 y2 0 x490 0 -0.182341597309204
Gyc2_491 y2 0 x491 0 0.113399279543516
Gyc2_492 y2 0 x492 0 0.0213667818340982
Gyc2_493 y2 0 x493 0 0.151313989015064
Gyc2_494 y2 0 x494 0 0.0587809424489495
Gyc2_495 y2 0 x495 0 0.0482749381940784
Gyc2_496 y2 0 x496 0 0.122773683416854
Gyc2_497 y2 0 x497 0 -0.0597955028291632
Gyc2_498 y2 0 x498 0 -0.0970976642155978
Gyc2_499 y2 0 x499 0 -0.0467974269720566
Gyc2_500 y2 0 x500 0 -0.0260208794876229
Gyc2_501 y2 0 x501 0 -0.214725530983838
Gyc2_502 y2 0 x502 0 -0.0284583880883695
Gyc2_503 y2 0 x503 0 -0.152221209250838
Gyc2_504 y2 0 x504 0 -0.361879684248225
Gyc2_505 y2 0 x505 0 -0.116705468007104
Gyc2_506 y2 0 x506 0 0.04441537000177
Gyc2_507 y2 0 x507 0 0.098598154495627
Gyc2_508 y2 0 x508 0 0.0661093952478097
Gyc2_509 y2 0 x509 0 0.22878164678056
Gyc2_510 y2 0 x510 0 -0.00992502462797449
Gyc2_511 y2 0 x511 0 -0.0965023255828883
Gyc2_512 y2 0 x512 0 -0.101091962875983
Gyc2_513 y2 0 x513 0 0.0821268790579624
Gyc2_514 y2 0 x514 0 -0.0686167855483267
Gyc2_515 y2 0 x515 0 -0.0391528824902644
Gyc2_516 y2 0 x516 0 -0.0320045378773161
Gyc2_517 y2 0 x517 0 -0.0921303480647536
Gyc2_518 y2 0 x518 0 -0.015553880211424
Gyc2_519 y2 0 x519 0 0.0733167203009233
Gyc2_520 y2 0 x520 0 -0.0150829867055327
Gyc2_521 y2 0 x521 0 0.0888578075042404
Gyc2_522 y2 0 x522 0 -0.0134269024007552
Gyc2_523 y2 0 x523 0 0.0568956792499786
Gyc2_524 y2 0 x524 0 -0.0518290080635309
Gyc2_525 y2 0 x525 0 0.0253931149123906
Gyc2_526 y2 0 x526 0 -0.0913254071352052
Gyc2_527 y2 0 x527 0 -0.0965891114469841
Gyc2_528 y2 0 x528 0 -0.0161716276489424
Gyc2_529 y2 0 x529 0 0.0898405063106121
Gyc2_530 y2 0 x530 0 0.017177223455059
Gyc2_531 y2 0 x531 0 -0.0783789181609506
Gyc2_532 y2 0 x532 0 0.0905112664639087
Gyc2_533 y2 0 x533 0 0.0862161510877341
Gyc2_534 y2 0 x534 0 0.0540072574154417
Gyc2_535 y2 0 x535 0 -0.112685557360637
Gyc2_536 y2 0 x536 0 0.120592671945346
Gyc2_537 y2 0 x537 0 -0.0667154903908046
Gyc2_538 y2 0 x538 0 0.104362499580185
Gyc2_539 y2 0 x539 0 0.0222704364578032
Gyc2_540 y2 0 x540 0 -0.120234215068773
Gyc2_541 y2 0 x541 0 -0.0229455491960522
Gyc2_542 y2 0 x542 0 0.0754175436389734
Gyc2_543 y2 0 x543 0 0.0878945681420245
Gyc2_544 y2 0 x544 0 0.221581424895071
Gyc2_545 y2 0 x545 0 -0.0610076077551971
Gyc2_546 y2 0 x546 0 -0.0253126844529137
Gyc2_547 y2 0 x547 0 -0.0399422940171444
Gyc2_548 y2 0 x548 0 1
Gyc2_549 y2 0 x549 0 0.0749346690957148
Gyc2_550 y2 0 x550 0 -0.0499363379048565
Gyc2_551 y2 0 x551 0 0.0737930435133163
Gyc2_552 y2 0 x552 0 -0.0888797227885077
Gyc2_553 y2 0 x553 0 0.0176764145161922
Gyc2_554 y2 0 x554 0 0.187085912060686
Gyc2_555 y2 0 x555 0 -0.0354601768939684
Gyc2_556 y2 0 x556 0 0.0392006611308457
Gyc2_557 y2 0 x557 0 -1
Gyc2_558 y2 0 x558 0 0.147148548421056
Gyc2_559 y2 0 x559 0 0.0333853817072219
Gyc2_560 y2 0 x560 0 -0.100740949269419
Gyc2_561 y2 0 x561 0 1
Gyc2_562 y2 0 x562 0 -0.0645140766960051
Gyc2_563 y2 0 x563 0 0.159093654492432
Gyc2_564 y2 0 x564 0 -0.0441578745212961
Gyc2_565 y2 0 x565 0 0.534443397285983
Gyc2_566 y2 0 x566 0 0.029834973083922
Gyc2_567 y2 0 x567 0 -0.092040348890806
Gyc2_568 y2 0 x568 0 -0.0420637163121097
Gyc2_569 y2 0 x569 0 -0.0859483534507027
Gyc2_570 y2 0 x570 0 0.0614611135966011
Gyc2_571 y2 0 x571 0 0.124588477159897
Gyc2_572 y2 0 x572 0 -0.0800008691873243
Gyc2_573 y2 0 x573 0 -0.924324333615379
Gyc2_574 y2 0 x574 0 0.0712602473500396
Gyc2_575 y2 0 x575 0 1
Gyc2_576 y2 0 x576 0 0.0586691994771216
Gyc2_577 y2 0 x577 0 0.102755662594436
Gyc2_578 y2 0 x578 0 -0.107563492581047
Gyc2_579 y2 0 x579 0 -0.107469674698705
Gyc2_580 y2 0 x580 0 0.0700297633050761
Gyc2_581 y2 0 x581 0 0.116793017254341
Gyc2_582 y2 0 x582 0 -0.00738952048269571
Gyc2_583 y2 0 x583 0 -0.332597350788244
Gyc2_584 y2 0 x584 0 -0.0446996234572574
Gyc2_585 y2 0 x585 0 -0.0390681318327677
Gyc2_586 y2 0 x586 0 -0.322774960775758
Gyc2_587 y2 0 x587 0 0.0926585852452756
Gyc2_588 y2 0 x588 0 0.111584883516874
Gyc2_589 y2 0 x589 0 -0.059063029052146
Gyc2_590 y2 0 x590 0 -0.109571780533375
Gyc2_591 y2 0 x591 0 0.0489670550745425
Gyc2_592 y2 0 x592 0 0.458578283881705
Gyc2_593 y2 0 x593 0 0.0868660256984451
Gyc2_594 y2 0 x594 0 -0.066086281799255
Gyc2_595 y2 0 x595 0 -0.087426208459677
Gyc2_596 y2 0 x596 0 -0.125359440775211
Gyc2_597 y2 0 x597 0 0.262686016441994
Gyc2_598 y2 0 x598 0 -0.147284304069315
Gyc2_599 y2 0 x599 0 0.0774886829733681
Gyc2_600 y2 0 x600 0 -0.146856903551446
Gyc2_601 y2 0 x601 0 -0.122338739658109
Gyc2_602 y2 0 x602 0 -0.00275151276629564
Gyc2_603 y2 0 x603 0 -0.203352404305611
Gyc2_604 y2 0 x604 0 0.109179987053025
Gyc2_605 y2 0 x605 0 0.107324527394449
Gyc2_606 y2 0 x606 0 -0.114857863212234
Gyc2_607 y2 0 x607 0 0.129856438038183
Gyc2_608 y2 0 x608 0 -0.0412370061854077
Gyc2_609 y2 0 x609 0 0.0677797946272793
Gyc2_610 y2 0 x610 0 0.0433920830879039
Gyc2_611 y2 0 x611 0 0.687172678463275
Gyc2_612 y2 0 x612 0 -0.094791023236451
Gyc2_613 y2 0 x613 0 -0.235302174927066
Gyc2_614 y2 0 x614 0 0.168335193227453
Gyc2_615 y2 0 x615 0 -0.315325366271665
Gyc2_616 y2 0 x616 0 -0.0130056720896154
Gyc2_617 y2 0 x617 0 -0.0189352211632178
Gyc2_618 y2 0 x618 0 0.15447662362207
Gyc2_619 y2 0 x619 0 -0.0907593350346678
Gyc2_620 y2 0 x620 0 0.0809451422853971
Gyc2_621 y2 0 x621 0 -0.105704826687975
Gyc2_622 y2 0 x622 0 0.109210444685561
Gyc2_623 y2 0 x623 0 0.418781024210194
Gyc2_624 y2 0 x624 0 -0.0621798343089405
Gyc2_625 y2 0 x625 0 0.0513315430140941
Gyc2_626 y2 0 x626 0 -0.0206193459348372
Gyc2_627 y2 0 x627 0 -0.0560486578855516
Gyc2_628 y2 0 x628 0 0.261152706032868
Gyc2_629 y2 0 x629 0 0.120093967870121
Gyc2_630 y2 0 x630 0 0.110553217880401
Gyc2_631 y2 0 x631 0 0.0840437496983336
Gyc2_632 y2 0 x632 0 -0.0244940454081787
Gyc2_633 y2 0 x633 0 0.0791710861050651
Gyc2_634 y2 0 x634 0 0.0894650444787266
Gyc2_635 y2 0 x635 0 -0.166302574342059
Gyc2_636 y2 0 x636 0 -0.104127221123196
Gyc2_637 y2 0 x637 0 0.0837596912212723
Gyc2_638 y2 0 x638 0 -0.0745664185590589
Gyc2_639 y2 0 x639 0 -0.0969104708608637
Gyc2_640 y2 0 x640 0 -0.0644530233028299
Gyc2_641 y2 0 x641 0 -0.17283088834303
Gyc2_642 y2 0 x642 0 0.0517392865986693
Gyc2_643 y2 0 x643 0 -0.0252144824275627
Gyc2_644 y2 0 x644 0 0.114930440224212
Gyc2_645 y2 0 x645 0 -0.0867428861087882
Gyc2_646 y2 0 x646 0 -0.0991291683226475
Gyc2_647 y2 0 x647 0 -0.106567182526592
Gyc2_648 y2 0 x648 0 -0.081162906123306
Gyc2_649 y2 0 x649 0 0.0967048061140728
Gyc2_650 y2 0 x650 0 -0.0601786897461999
Gyc2_651 y2 0 x651 0 -0.0898733849289913
Gyc2_652 y2 0 x652 0 -0.141662629510802
Gyc2_653 y2 0 x653 0 -0.0568221071908808
Gyc2_654 y2 0 x654 0 -0.07495904166114
Gyc2_655 y2 0 x655 0 -0.315146907201803
Gyc2_656 y2 0 x656 0 0.253702105757671
Gyc2_657 y2 0 x657 0 -0.101313082361356
Gyc2_658 y2 0 x658 0 -0.0843848047599242
Gyc2_659 y2 0 x659 0 -0.000656219164256508
Gyc2_660 y2 0 x660 0 0.0678396971363599
Gyc2_661 y2 0 x661 0 -0.16939919901724
Gyc2_662 y2 0 x662 0 0.0998163073681342
Gyc2_663 y2 0 x663 0 0.0262091139641673
Gyc2_664 y2 0 x664 0 -0.118622374639814
Gyc2_665 y2 0 x665 0 0.0439915795951888
Gyc2_666 y2 0 x666 0 -0.0108364864555495
Gyc2_667 y2 0 x667 0 -0.0480164370868879
Gyc2_668 y2 0 x668 0 0.125661267360811
Gyc2_669 y2 0 x669 0 -0.0774894073905441
Gyc2_670 y2 0 x670 0 -0.1041102937563
Gyc2_671 y2 0 x671 0 -0.148672243085698
Gyc2_672 y2 0 x672 0 0.123870571811127
Gyc2_673 y2 0 x673 0 -0.0805585213880285
Gyc2_674 y2 0 x674 0 -0.110428263891053
Gyc2_675 y2 0 x675 0 0.0708872227540954
Gyc2_676 y2 0 x676 0 0.109429494932908
Gyc2_677 y2 0 x677 0 0.0409988645612391
Gyc2_678 y2 0 x678 0 -0.0510779824450801
Gyc2_679 y2 0 x679 0 0.0850016288708968
Gyc2_680 y2 0 x680 0 -0.0873867331145546
Gyc2_681 y2 0 x681 0 0.0515700352287419
Gyc2_682 y2 0 x682 0 -0.10407346257317
Gyc2_683 y2 0 x683 0 -0.0912927033997605
Gyc2_684 y2 0 x684 0 0.00827304686210106
Gyc2_685 y2 0 x685 0 0.119679955057338
Gyc2_686 y2 0 x686 0 0.110619479657292
Gyc2_687 y2 0 x687 0 0.0484602679397039
Gyc2_688 y2 0 x688 0 -0.0992329646827662
Gyc2_689 y2 0 x689 0 0.0974128912659078
Gyc2_690 y2 0 x690 0 -1
Gyc2_691 y2 0 x691 0 0.107004155937082
Gyc2_692 y2 0 x692 0 -0.0971970894198887
Gyc2_693 y2 0 x693 0 0.100812390645135
Gyc2_694 y2 0 x694 0 0.242419609436653
Gyc2_695 y2 0 x695 0 -0.069697432371335
Gyc2_696 y2 0 x696 0 0.118041617489206
Gyc2_697 y2 0 x697 0 -0.0644123054890555
Gyc2_698 y2 0 x698 0 -0.0303415376886174
Gyc2_699 y2 0 x699 0 -1
Gyc2_700 y2 0 x700 0 0.03546431813454
Gyc2_701 y2 0 x701 0 0.127958643077578
Gyc2_702 y2 0 x702 0 0.124323586212416
Gyc2_703 y2 0 x703 0 -0.235142963887532
Gyc2_704 y2 0 x704 0 -0.120554049447538
Gyc2_705 y2 0 x705 0 -0.109272747980753
Gyc2_706 y2 0 x706 0 0.12023066343991
Gyc2_707 y2 0 x707 0 -0.133424199179449
Gyc2_708 y2 0 x708 0 0.11903240646541
Gyc2_709 y2 0 x709 0 -0.143084885064205
Gyc2_710 y2 0 x710 0 0.216525145985962
Gyc2_711 y2 0 x711 0 0.0292695476396624
Gyc2_712 y2 0 x712 0 -0.166530977340039
Gyc2_713 y2 0 x713 0 -0.114141035920484
Gyc2_714 y2 0 x714 0 1
Gyc2_715 y2 0 x715 0 -0.103173480540368
Gyc2_716 y2 0 x716 0 0.0810856267050483
Gyc2_717 y2 0 x717 0 0.0843091773310129
Gyc2_718 y2 0 x718 0 -0.0993397968638064
Gyc2_719 y2 0 x719 0 -0.0826469257396643
Gyc2_720 y2 0 x720 0 0.0834011679137504
Gyc2_721 y2 0 x721 0 0.252411176956799
Gyc2_722 y2 0 x722 0 0.0590663743205447
Gyc2_723 y2 0 x723 0 -0.0220938104497508
Gyc2_724 y2 0 x724 0 -0.00118062325779979
Gyc2_725 y2 0 x725 0 -0.0987673375428721
Gyc2_726 y2 0 x726 0 0.0219292722130962
Gyc2_727 y2 0 x727 0 0.199405454902599
Gyc2_728 y2 0 x728 0 0.012768110283363
Gyc2_729 y2 0 x729 0 -0.0912827077193226
Gyc2_730 y2 0 x730 0 0.105299861644167
Gyc2_731 y2 0 x731 0 -0.0860520653393504
Gyc2_732 y2 0 x732 0 0.0989048856528331
Gyc2_733 y2 0 x733 0 0.121366807754154
Gyc2_734 y2 0 x734 0 0.0925317625520899
Gyc2_735 y2 0 x735 0 -1
Gyc2_736 y2 0 x736 0 -0.075162999595538
Gyc2_737 y2 0 x737 0 0.104323975310536
Gyc2_738 y2 0 x738 0 0.0247634735219906
Gyc2_739 y2 0 x739 0 0.0977695830676691
Gyc2_740 y2 0 x740 0 0.0955660301158605
Gyc2_741 y2 0 x741 0 -0.745542364966214
Gyc2_742 y2 0 x742 0 -0.0702845522277359
Gyc2_743 y2 0 x743 0 -0.0155938798242585
Gyc2_744 y2 0 x744 0 0.104595556282403
Gyc2_745 y2 0 x745 0 -0.0918967916674041
Gyc2_746 y2 0 x746 0 -0.16672911467857
Gyc2_747 y2 0 x747 0 -0.0564813557051069
Gyc2_748 y2 0 x748 0 1
Gyc2_749 y2 0 x749 0 -0.0985286046625027
Gyc2_750 y2 0 x750 0 0.598238667297851
Gyc2_751 y2 0 x751 0 -0.0931766056168719
Gyc2_752 y2 0 x752 0 -0.0857729392357868
Gyc2_753 y2 0 x753 0 -0.0656665143495242
Gyc2_754 y2 0 x754 0 0.11638158575697
Gyc2_755 y2 0 x755 0 0.114326091648084
Gyc2_756 y2 0 x756 0 -0.099132506989164
Gyc2_757 y2 0 x757 0 0.125599013256546
Gyc2_758 y2 0 x758 0 0.0940737303650728
Gyc2_759 y2 0 x759 0 0.0616836246361804
Gyc2_760 y2 0 x760 0 -0.278169811771896
Gyc2_761 y2 0 x761 0 0.108040484948898
Gyc2_762 y2 0 x762 0 -0.0864720662896779
Gyc2_763 y2 0 x763 0 -0.101950931379713
Gyc2_764 y2 0 x764 0 -0.0955317437032919
Gyc2_765 y2 0 x765 0 0.0588954778781226
Gyc2_766 y2 0 x766 0 -0.0255641260011063
Gyc2_767 y2 0 x767 0 -0.116846490760146
Gyc2_768 y2 0 x768 0 0.078125054178974
Gyc2_769 y2 0 x769 0 0.0782737390662519
Gyc2_770 y2 0 x770 0 -0.0815560946343585
Gyc2_771 y2 0 x771 0 0.107186477076964
Gyc2_772 y2 0 x772 0 0.0964561913862441
Gyc2_773 y2 0 x773 0 0.115864842494277
Gyc2_774 y2 0 x774 0 0.167353393762982
Gyc2_775 y2 0 x775 0 0.447228937671219
Gyc2_776 y2 0 x776 0 0.152741149049744
Gyc2_777 y2 0 x777 0 -0.0625718183964559
Gyc2_778 y2 0 x778 0 0.112520569816898
Gyc2_779 y2 0 x779 0 0.0909600656261173
Gyc2_780 y2 0 x780 0 0.76487290126911
Gyc2_781 y2 0 x781 0 0.0709152016012379
Gyc2_782 y2 0 x782 0 0.10245890426368
Gyc2_783 y2 0 x783 0 0.0974576139279935
Gyc2_784 y2 0 x784 0 -0.0428373775711032
Gyc2_785 y2 0 x785 0 0.114921483972856
Gyc2_786 y2 0 x786 0 -0.0963086745665744
Gyc2_787 y2 0 x787 0 -0.0555348293386092
Gyc2_788 y2 0 x788 0 -0.0845940309825825
Gyc2_789 y2 0 x789 0 -0.113623838619616
Gyc2_790 y2 0 x790 0 0.733592224692746
Gyc2_791 y2 0 x791 0 -0.0704779655715486
Gyc2_792 y2 0 x792 0 -0.107304020197839
Gyc2_793 y2 0 x793 0 0.2437699430779
Gyc2_794 y2 0 x794 0 0.162762768793503
Gyc2_795 y2 0 x795 0 -0.0915045918764373
Gyc2_796 y2 0 x796 0 -0.0874775279068651
Gyc2_797 y2 0 x797 0 0.0108480065180583
Gyc2_798 y2 0 x798 0 0.0435108608790306
Gyc2_799 y2 0 x799 0 -0.0766334757177766
Gyc2_800 y2 0 x800 0 0.0802832638844148
Gyc2_801 y2 0 x801 0 -0.777480190818726
Gyc2_802 y2 0 x802 0 -1
Gyc2_803 y2 0 x803 0 1
Gyc2_804 y2 0 x804 0 -1
Gyc2_805 y2 0 x805 0 -1
Gyc2_806 y2 0 x806 0 -1
Gyc2_807 y2 0 x807 0 1
Gyc2_808 y2 0 x808 0 1
Gyc2_809 y2 0 x809 0 -1
Gyc2_810 y2 0 x810 0 1
Gyc2_811 y2 0 x811 0 1
Gyc2_812 y2 0 x812 0 1
Gyc2_813 y2 0 x813 0 1
Gyc2_814 y2 0 x814 0 -1
Gyc2_815 y2 0 x815 0 1
Gyc2_816 y2 0 x816 0 1
Gyc2_817 y2 0 x817 0 1
Gyc2_818 y2 0 x818 0 -1
Gyc2_819 y2 0 x819 0 1
Gyc2_820 y2 0 x820 0 1
Gyc2_821 y2 0 x821 0 1
Gyc2_822 y2 0 x822 0 -1
Gyc2_823 y2 0 x823 0 -1
Gyc2_824 y2 0 x824 0 -1
Gyc2_825 y2 0 x825 0 -1
Gyc2_826 y2 0 x826 0 -1
Gyc2_827 y2 0 x827 0 1
Gyc2_828 y2 0 x828 0 -1
Gyc2_829 y2 0 x829 0 1
Gyc2_830 y2 0 x830 0 -1
Gyc2_831 y2 0 x831 0 1
Gyc2_832 y2 0 x832 0 -1
Gyc2_833 y2 0 x833 0 1
Gyc2_834 y2 0 x834 0 -1
Gyc2_835 y2 0 x835 0 1
Gyc2_836 y2 0 x836 0 -1
Gyc2_837 y2 0 x837 0 -1
Gyc2_838 y2 0 x838 0 1
Gyc2_839 y2 0 x839 0 -1
Gyc2_840 y2 0 x840 0 1
Gyc2_841 y2 0 x841 0 1
Gyc2_842 y2 0 x842 0 -1
Gyc2_843 y2 0 x843 0 1
Gyc2_844 y2 0 x844 0 1
Gyc2_845 y2 0 x845 0 1
Gyc2_846 y2 0 x846 0 -1
Gyc2_847 y2 0 x847 0 1
Gyc2_848 y2 0 x848 0 -1
Gyc2_849 y2 0 x849 0 -1
Gyc2_850 y2 0 x850 0 -1
Gyc2_851 y2 0 x851 0 1
Gyc2_852 y2 0 x852 0 1
Gyc2_853 y2 0 x853 0 1
Gyc2_854 y2 0 x854 0 -1
Gyc2_855 y2 0 x855 0 1
Gyc2_856 y2 0 x856 0 -1
Gyc2_857 y2 0 x857 0 1
Gyc2_858 y2 0 x858 0 1
Gyc2_859 y2 0 x859 0 -1
Gyc2_860 y2 0 x860 0 -1
Gyc2_861 y2 0 x861 0 -1
Gyc2_862 y2 0 x862 0 1
Gyc2_863 y2 0 x863 0 -1
Gyc2_864 y2 0 x864 0 1
Gyc2_865 y2 0 x865 0 1
Gyc2_866 y2 0 x866 0 1
Gyc2_867 y2 0 x867 0 1
Gyc2_868 y2 0 x868 0 -1
Gyc2_869 y2 0 x869 0 1
Gyc2_870 y2 0 x870 0 -1
Gyc2_871 y2 0 x871 0 -1
Gyc2_872 y2 0 x872 0 1
Gyc2_873 y2 0 x873 0 -1
Gyc2_874 y2 0 x874 0 1
Gyc2_875 y2 0 x875 0 -1
Gyc2_876 y2 0 x876 0 -1
Gyc2_877 y2 0 x877 0 -1
Gyc2_878 y2 0 x878 0 1
Gyc2_879 y2 0 x879 0 1
Gyc2_880 y2 0 x880 0 -1
Gyc2_881 y2 0 x881 0 1
Gyc2_882 y2 0 x882 0 1
Gyc2_883 y2 0 x883 0 -1
Gyc2_884 y2 0 x884 0 1
Gyc2_885 y2 0 x885 0 -1
Gyc2_886 y2 0 x886 0 1
Gyc2_887 y2 0 x887 0 1
Gyc2_888 y2 0 x888 0 1
Gyc2_889 y2 0 x889 0 -1
Gyc2_890 y2 0 x890 0 1
Gyc2_891 y2 0 x891 0 1
Gyc2_892 y2 0 x892 0 1
Gyc2_893 y2 0 x893 0 -0.00123198099303243
Gyc2_894 y2 0 x894 0 1
Gyc2_895 y2 0 x895 0 -1
Gyc2_896 y2 0 x896 0 -1
Gyc2_897 y2 0 x897 0 -1
Gyc2_898 y2 0 x898 0 -1
Gyc2_899 y2 0 x899 0 -1
Gyc2_900 y2 0 x900 0 -1
Gyc2_901 y2 0 x901 0 -0.503827114401445
Gyc2_902 y2 0 x902 0 -1
Gyc2_903 y2 0 x903 0 -1
Gyc2_904 y2 0 x904 0 -1
Gyc2_905 y2 0 x905 0 -1
Gyc2_906 y2 0 x906 0 1
Gyc2_907 y2 0 x907 0 -1
Gyc2_908 y2 0 x908 0 1
Gyc2_909 y2 0 x909 0 -1
Gyc2_910 y2 0 x910 0 -1
Gyc2_911 y2 0 x911 0 -1
Gyc2_912 y2 0 x912 0 1
Gyc2_913 y2 0 x913 0 -1
Gyc2_914 y2 0 x914 0 1
Gyc2_915 y2 0 x915 0 -1
Gyc2_916 y2 0 x916 0 1
Gyc2_917 y2 0 x917 0 1
Gyc2_918 y2 0 x918 0 1
Gyc2_919 y2 0 x919 0 1
Gyc2_920 y2 0 x920 0 1
Gyc2_921 y2 0 x921 0 1
Gyc2_922 y2 0 x922 0 -1
Gyc2_923 y2 0 x923 0 -1
Gyc2_924 y2 0 x924 0 -1
Gyc2_925 y2 0 x925 0 1
Gyc2_926 y2 0 x926 0 -1
Gyc2_927 y2 0 x927 0 -1
Gyc2_928 y2 0 x928 0 -1
Gyc2_929 y2 0 x929 0 -1
Gyc2_930 y2 0 x930 0 -1
Gyc2_931 y2 0 x931 0 1
Gyc2_932 y2 0 x932 0 -1
Gyc2_933 y2 0 x933 0 1
Gyc2_934 y2 0 x934 0 1
Gyc2_935 y2 0 x935 0 -1
Gyc2_936 y2 0 x936 0 -1
Gyc2_937 y2 0 x937 0 -1
Gyc2_938 y2 0 x938 0 1
Gyc2_939 y2 0 x939 0 -1
Gyc2_940 y2 0 x940 0 1
Gyc2_941 y2 0 x941 0 1
Gyc2_942 y2 0 x942 0 -1
Gyc2_943 y2 0 x943 0 -1
Gyc2_944 y2 0 x944 0 -1
Gyc2_945 y2 0 x945 0 1
Gyc2_946 y2 0 x946 0 1
Gyc2_947 y2 0 x947 0 1
Gyc2_948 y2 0 x948 0 1
Gyc2_949 y2 0 x949 0 1
Gyc2_950 y2 0 x950 0 -1
Gyc2_951 y2 0 x951 0 -1
Gyc2_952 y2 0 x952 0 -1
Gyc2_953 y2 0 x953 0 1
Gyc2_954 y2 0 x954 0 -1
Gyc2_955 y2 0 x955 0 1
Gyc2_956 y2 0 x956 0 1
Gyc2_957 y2 0 x957 0 1
Gyc2_958 y2 0 x958 0 1
Gyc2_959 y2 0 x959 0 -1
Gyc2_960 y2 0 x960 0 1
Gyc2_961 y2 0 x961 0 1
Gyc2_962 y2 0 x962 0 -1
Gyc2_963 y2 0 x963 0 1
Gyc2_964 y2 0 x964 0 -1
Gyc2_965 y2 0 x965 0 -1
Gyc2_966 y2 0 x966 0 1
Gyc2_967 y2 0 x967 0 -1
Gyc2_968 y2 0 x968 0 -1
Gyc2_969 y2 0 x969 0 1
Gyc2_970 y2 0 x970 0 1
Gyc2_971 y2 0 x971 0 -1
Gyc2_972 y2 0 x972 0 1
Gyc2_973 y2 0 x973 0 1
Gyc2_974 y2 0 x974 0 -1
Gyc2_975 y2 0 x975 0 -1
Gyc2_976 y2 0 x976 0 1
Gyc2_977 y2 0 x977 0 1
Gyc2_978 y2 0 x978 0 -1
Gyc2_979 y2 0 x979 0 1
Gyc2_980 y2 0 x980 0 1
Gyc2_981 y2 0 x981 0 -1
Gyc2_982 y2 0 x982 0 -1
Gyc2_983 y2 0 x983 0 -1
Gyc2_984 y2 0 x984 0 1
Gyc2_985 y2 0 x985 0 -1
Gyc2_986 y2 0 x986 0 1
Gyc2_987 y2 0 x987 0 -1
Gyc2_988 y2 0 x988 0 -1
Gyc2_989 y2 0 x989 0 -1
Gyc2_990 y2 0 x990 0 -1
Gyc2_991 y2 0 x991 0 -1
Gyc2_992 y2 0 x992 0 -1
Gyc2_993 y2 0 x993 0 -1
Gyc2_994 y2 0 x994 0 1
Gyc2_995 y2 0 x995 0 1
Gyc2_996 y2 0 x996 0 1
Gyc2_997 y2 0 x997 0 -1
Gyc2_998 y2 0 x998 0 -1
Gyc2_999 y2 0 x999 0 -1
Gyc2_1000 y2 0 x1000 0 -1
Gyc2_1001 y2 0 x1001 0 -1
Gyc2_1002 y2 0 x1002 0 -1
Gyc2_1003 y2 0 x1003 0 1
Gyc2_1004 y2 0 x1004 0 -1
Gyc2_1005 y2 0 x1005 0 1
Gyc2_1006 y2 0 x1006 0 -1
Gyc2_1007 y2 0 x1007 0 -1
Gyc2_1008 y2 0 x1008 0 1
Gyc2_1009 y2 0 x1009 0 1
Gyc2_1010 y2 0 x1010 0 -1
Gyc2_1011 y2 0 x1011 0 -1
Gyc2_1012 y2 0 x1012 0 1
Gyc2_1013 y2 0 x1013 0 -1
Gyc2_1014 y2 0 x1014 0 -1
Gyc2_1015 y2 0 x1015 0 -1
Gyc2_1016 y2 0 x1016 0 -1
Gyc2_1017 y2 0 x1017 0 1
Gyc2_1018 y2 0 x1018 0 -1
Gyc2_1019 y2 0 x1019 0 -1
Gyc2_1020 y2 0 x1020 0 -1
Gyc2_1021 y2 0 x1021 0 1
Gyc2_1022 y2 0 x1022 0 1
Gyc2_1023 y2 0 x1023 0 -1
Gyc2_1024 y2 0 x1024 0 1
Gyc2_1025 y2 0 x1025 0 -1
Gyc2_1026 y2 0 x1026 0 1
Gyc2_1027 y2 0 x1027 0 -1
Gyc2_1028 y2 0 x1028 0 1
Gyc2_1029 y2 0 x1029 0 -1
Gyc2_1030 y2 0 x1030 0 1
Gyc2_1031 y2 0 x1031 0 1
Gyc2_1032 y2 0 x1032 0 1
Gyc2_1033 y2 0 x1033 0 1
Gyc2_1034 y2 0 x1034 0 1
Gyc2_1035 y2 0 x1035 0 1
Gyc2_1036 y2 0 x1036 0 -1
Gyc2_1037 y2 0 x1037 0 -1
Gyc2_1038 y2 0 x1038 0 -1
Gyc2_1039 y2 0 x1039 0 -0.0941717777321933
Gyc2_1040 y2 0 x1040 0 -1
Gyc2_1041 y2 0 x1041 0 -1
Gyc2_1042 y2 0 x1042 0 -1
Gyc2_1043 y2 0 x1043 0 1
Gyc2_1044 y2 0 x1044 0 -1
Gyc2_1045 y2 0 x1045 0 1
Gyc2_1046 y2 0 x1046 0 1
Gyc2_1047 y2 0 x1047 0 -1
Gyc2_1048 y2 0 x1048 0 1
Gyc2_1049 y2 0 x1049 0 1
Gyc2_1050 y2 0 x1050 0 -1
Gyc2_1051 y2 0 x1051 0 -1
Gyc2_1052 y2 0 x1052 0 -1
Gyc2_1053 y2 0 x1053 0 1
Gyc2_1054 y2 0 x1054 0 -1
Gyc2_1055 y2 0 x1055 0 -1
Gyc2_1056 y2 0 x1056 0 1
Gyc2_1057 y2 0 x1057 0 -1
Gyc2_1058 y2 0 x1058 0 -1
Gyc2_1059 y2 0 x1059 0 -1
Gyc2_1060 y2 0 x1060 0 1
Gyc2_1061 y2 0 x1061 0 -1
Gyc2_1062 y2 0 x1062 0 1
Gyc2_1063 y2 0 x1063 0 1
Gyc2_1064 y2 0 x1064 0 1
Gyc2_1065 y2 0 x1065 0 -1
Gyc2_1066 y2 0 x1066 0 -1
Gyc2_1067 y2 0 x1067 0 -1
Gyc2_1068 y2 0 x1068 0 -1
Gyc2_1069 y2 0 x1069 0 1
Gyc2_1070 y2 0 x1070 0 -1
Gyc2_1071 y2 0 x1071 0 1
Gyc2_1072 y2 0 x1072 0 1
Gyc2_1073 y2 0 x1073 0 1
Gyc2_1074 y2 0 x1074 0 -1
Gyc2_1075 y2 0 x1075 0 1
Gyc2_1076 y2 0 x1076 0 -1
Gyc2_1077 y2 0 x1077 0 -1
Gyc2_1078 y2 0 x1078 0 -1
Gyc2_1079 y2 0 x1079 0 -1
Gyc2_1080 y2 0 x1080 0 -1
Gyc2_1081 y2 0 x1081 0 1
Gyc2_1082 y2 0 x1082 0 1
Gyc2_1083 y2 0 x1083 0 -1
Gyc2_1084 y2 0 x1084 0 1
Gyc2_1085 y2 0 x1085 0 -1
Gyc2_1086 y2 0 x1086 0 1
Gyc2_1087 y2 0 x1087 0 -1
Gyc2_1088 y2 0 x1088 0 -1
Gyc2_1089 y2 0 x1089 0 -1
Gyc2_1090 y2 0 x1090 0 -1
Gyc2_1091 y2 0 x1091 0 1
Gyc2_1092 y2 0 x1092 0 1
Gyc2_1093 y2 0 x1093 0 1
Gyc2_1094 y2 0 x1094 0 1
Gyc2_1095 y2 0 x1095 0 1
Gyc2_1096 y2 0 x1096 0 -1
Gyc2_1097 y2 0 x1097 0 1
Gyc2_1098 y2 0 x1098 0 -1
Gyc2_1099 y2 0 x1099 0 1
Gyc2_1100 y2 0 x1100 0 -1
Gyc2_1101 y2 0 x1101 0 -1
Gyc2_1102 y2 0 x1102 0 -1
Gyc2_1103 y2 0 x1103 0 -1
Gyc2_1104 y2 0 x1104 0 1
Gyc2_1105 y2 0 x1105 0 1
Gyc2_1106 y2 0 x1106 0 1
Gyc2_1107 y2 0 x1107 0 1
Gyc2_1108 y2 0 x1108 0 1
Gyc2_1109 y2 0 x1109 0 -1
Gyc2_1110 y2 0 x1110 0 -1
Gyc2_1111 y2 0 x1111 0 -1
Gyc2_1112 y2 0 x1112 0 -1
Gyc2_1113 y2 0 x1113 0 1
Gyc2_1114 y2 0 x1114 0 -1
Gyc2_1115 y2 0 x1115 0 1
Gyc2_1116 y2 0 x1116 0 1
Gyc2_1117 y2 0 x1117 0 1
Gyc2_1118 y2 0 x1118 0 -1
Gyc2_1119 y2 0 x1119 0 1
Gyc2_1120 y2 0 x1120 0 -1
Gyc2_1121 y2 0 x1121 0 1
Gyc2_1122 y2 0 x1122 0 1
Gyc2_1123 y2 0 x1123 0 1
Gyc2_1124 y2 0 x1124 0 1
Gyc2_1125 y2 0 x1125 0 -1
Gyc2_1126 y2 0 x1126 0 -1
Gyc2_1127 y2 0 x1127 0 1
Gyc2_1128 y2 0 x1128 0 1
Gyc2_1129 y2 0 x1129 0 1
Gyc2_1130 y2 0 x1130 0 1
Gyc2_1131 y2 0 x1131 0 1
Gyc2_1132 y2 0 x1132 0 1
Gyc2_1133 y2 0 x1133 0 1
Gyc2_1134 y2 0 x1134 0 1
Gyc2_1135 y2 0 x1135 0 1
Gyc2_1136 y2 0 x1136 0 1
Gyc2_1137 y2 0 x1137 0 1
Gyc2_1138 y2 0 x1138 0 -1
Gyc2_1139 y2 0 x1139 0 1
Gyc2_1140 y2 0 x1140 0 -1
Gyc2_1141 y2 0 x1141 0 -1
Gyc2_1142 y2 0 x1142 0 -1
Gyc2_1143 y2 0 x1143 0 1
Gyc2_1144 y2 0 x1144 0 1
Gyc2_1145 y2 0 x1145 0 1
Gyc2_1146 y2 0 x1146 0 1
Gyc2_1147 y2 0 x1147 0 1
Gyc2_1148 y2 0 x1148 0 -1
Gyc2_1149 y2 0 x1149 0 1
Gyc2_1150 y2 0 x1150 0 1
Gyc2_1151 y2 0 x1151 0 1
Gyc2_1152 y2 0 x1152 0 -1
Gyc2_1153 y2 0 x1153 0 -1
Gyc2_1154 y2 0 x1154 0 1
Gyc2_1155 y2 0 x1155 0 1
Gyc2_1156 y2 0 x1156 0 -1
Gyc2_1157 y2 0 x1157 0 -1
Gyc2_1158 y2 0 x1158 0 -1
Gyc2_1159 y2 0 x1159 0 -1
Gyc2_1160 y2 0 x1160 0 -1
Gyc2_1161 y2 0 x1161 0 1
Gyc2_1162 y2 0 x1162 0 -1
Gyc2_1163 y2 0 x1163 0 1
Gyc2_1164 y2 0 x1164 0 -1
Gyc2_1165 y2 0 x1165 0 1
Gyc2_1166 y2 0 x1166 0 1
Gyc2_1167 y2 0 x1167 0 1
Gyc2_1168 y2 0 x1168 0 -1
Gyc2_1169 y2 0 x1169 0 -1
Gyc2_1170 y2 0 x1170 0 -1
Gyc2_1171 y2 0 x1171 0 -1
Gyc2_1172 y2 0 x1172 0 1
Gyc2_1173 y2 0 x1173 0 1
Gyc2_1174 y2 0 x1174 0 1
Gyc2_1175 y2 0 x1175 0 1
Gyc2_1176 y2 0 x1176 0 1
Gyc2_1177 y2 0 x1177 0 1
Gyc2_1178 y2 0 x1178 0 -1
Gyc2_1179 y2 0 x1179 0 1
Gyc2_1180 y2 0 x1180 0 -1
Gyc2_1181 y2 0 x1181 0 -1
Gyc2_1182 y2 0 x1182 0 1
Gyc2_1183 y2 0 x1183 0 -1
Gyc2_1184 y2 0 x1184 0 1
Gyc2_1185 y2 0 x1185 0 -1
Gyc2_1186 y2 0 x1186 0 -1
Gyc2_1187 y2 0 x1187 0 1
Gyc2_1188 y2 0 x1188 0 -1
Gyc2_1189 y2 0 x1189 0 -1
Gyc2_1190 y2 0 x1190 0 -1
Gyc2_1191 y2 0 x1191 0 -1
Gyc2_1192 y2 0 x1192 0 1
Gyc2_1193 y2 0 x1193 0 -1
Gyc2_1194 y2 0 x1194 0 -1
Gyc2_1195 y2 0 x1195 0 -1
Gyc2_1196 y2 0 x1196 0 1
Gyc2_1197 y2 0 x1197 0 1
Gyc2_1198 y2 0 x1198 0 -1
Gyc2_1199 y2 0 x1199 0 -1
Gyc2_1200 y2 0 x1200 0 -1
Gyc2_1201 y2 0 x1201 0 1
Gyc2_1202 y2 0 x1202 0 1
Gyc2_1203 y2 0 x1203 0 -1
Gyc2_1204 y2 0 x1204 0 1
Gyc2_1205 y2 0 x1205 0 -1
Gyc2_1206 y2 0 x1206 0 1
Gyc2_1207 y2 0 x1207 0 1
Gyc2_1208 y2 0 x1208 0 -1
Gyc2_1209 y2 0 x1209 0 1
Gyc2_1210 y2 0 x1210 0 1
Gyc2_1211 y2 0 x1211 0 1
Gyc2_1212 y2 0 x1212 0 1
Gyc2_1213 y2 0 x1213 0 1
Gyc2_1214 y2 0 x1214 0 1
Gyc2_1215 y2 0 x1215 0 -1
Gyc2_1216 y2 0 x1216 0 1
Gyc2_1217 y2 0 x1217 0 1
Gyc2_1218 y2 0 x1218 0 -1
Gyc2_1219 y2 0 x1219 0 -1
Gyc2_1220 y2 0 x1220 0 -1
Gyc2_1221 y2 0 x1221 0 -1
Gyc2_1222 y2 0 x1222 0 1
Gyc2_1223 y2 0 x1223 0 1
Gyc2_1224 y2 0 x1224 0 -1
Gyc2_1225 y2 0 x1225 0 -1
Gyc2_1226 y2 0 x1226 0 1
Gyc2_1227 y2 0 x1227 0 -1
Gyc2_1228 y2 0 x1228 0 1
Gyc2_1229 y2 0 x1229 0 -1
Gyc2_1230 y2 0 x1230 0 1
Gyc2_1231 y2 0 x1231 0 -1
Gyc2_1232 y2 0 x1232 0 -1
Gyc2_1233 y2 0 x1233 0 -1
Gyc2_1234 y2 0 x1234 0 1
Gyc2_1235 y2 0 x1235 0 -1
Gyc2_1236 y2 0 x1236 0 1
Gyc2_1237 y2 0 x1237 0 1
Gyc2_1238 y2 0 x1238 0 -1
Gyc2_1239 y2 0 x1239 0 1
Gyc2_1240 y2 0 x1240 0 1
Gyc2_1241 y2 0 x1241 0 -1
Gyc2_1242 y2 0 x1242 0 1
Gyc2_1243 y2 0 x1243 0 1
Gyc2_1244 y2 0 x1244 0 -1
Gyc2_1245 y2 0 x1245 0 -1
Gyc2_1246 y2 0 x1246 0 -1
Gyc2_1247 y2 0 x1247 0 -1
Gyc2_1248 y2 0 x1248 0 1
Gyc2_1249 y2 0 x1249 0 1
Gyc2_1250 y2 0 x1250 0 -1
Gyc2_1251 y2 0 x1251 0 1
Gyc2_1252 y2 0 x1252 0 1
Gyc2_1253 y2 0 x1253 0 1
Gyc2_1254 y2 0 x1254 0 -1
Gyc2_1255 y2 0 x1255 0 1
Gyc2_1256 y2 0 x1256 0 -1
Gyc2_1257 y2 0 x1257 0 -1
Gyc2_1258 y2 0 x1258 0 1
Gyc2_1259 y2 0 x1259 0 -1
Gyc2_1260 y2 0 x1260 0 -1
Gyc2_1261 y2 0 x1261 0 -1
Gyc2_1262 y2 0 x1262 0 1
Gyc2_1263 y2 0 x1263 0 -1
Gyc2_1264 y2 0 x1264 0 1
Gyc2_1265 y2 0 x1265 0 1
Gyc2_1266 y2 0 x1266 0 1
Gyc2_1267 y2 0 x1267 0 1
Gyc2_1268 y2 0 x1268 0 -1
Gyc2_1269 y2 0 x1269 0 1
Gyc2_1270 y2 0 x1270 0 -1
Gyc2_1271 y2 0 x1271 0 1
Gyc2_1272 y2 0 x1272 0 -1
Gyc2_1273 y2 0 x1273 0 -1
Gyc2_1274 y2 0 x1274 0 1
Gyc2_1275 y2 0 x1275 0 -1
Gyc2_1276 y2 0 x1276 0 1
Gyc2_1277 y2 0 x1277 0 -1
Gyc2_1278 y2 0 x1278 0 1
Gyc2_1279 y2 0 x1279 0 -1
Gyc2_1280 y2 0 x1280 0 -1
Gyc2_1281 y2 0 x1281 0 -1
Gyc2_1282 y2 0 x1282 0 1
Gyc2_1283 y2 0 x1283 0 -1
Gyc2_1284 y2 0 x1284 0 1
Gyc2_1285 y2 0 x1285 0 1
Gyc2_1286 y2 0 x1286 0 -1
Gyc2_1287 y2 0 x1287 0 1
Gyc2_1288 y2 0 x1288 0 -1
Gyc2_1289 y2 0 x1289 0 -1
Gyc2_1290 y2 0 x1290 0 1
Gyc2_1291 y2 0 x1291 0 -1
Gyc2_1292 y2 0 x1292 0 1
Gyc2_1293 y2 0 x1293 0 -1
Gyc2_1294 y2 0 x1294 0 1
Gyc2_1295 y2 0 x1295 0 1
Gyc2_1296 y2 0 x1296 0 1
Gyc2_1297 y2 0 x1297 0 1
Gyc2_1298 y2 0 x1298 0 -1
Gyc2_1299 y2 0 x1299 0 -1
Gyc2_1300 y2 0 x1300 0 1
Gyc2_1301 y2 0 x1301 0 -1
Gyc2_1302 y2 0 x1302 0 1
Gyc2_1303 y2 0 x1303 0 -1
Gyc2_1304 y2 0 x1304 0 -1
Gyc2_1305 y2 0 x1305 0 -1
Gyc2_1306 y2 0 x1306 0 -1
Gyc2_1307 y2 0 x1307 0 1
Gyc2_1308 y2 0 x1308 0 1
Gyc2_1309 y2 0 x1309 0 1
Gyc2_1310 y2 0 x1310 0 1
Gyc2_1311 y2 0 x1311 0 -1
Gyc2_1312 y2 0 x1312 0 -1
Gyc2_1313 y2 0 x1313 0 -1
Gyc2_1314 y2 0 x1314 0 1
Gyc2_1315 y2 0 x1315 0 -1
Gyc2_1316 y2 0 x1316 0 1
Gyc2_1317 y2 0 x1317 0 -1
Gyc2_1318 y2 0 x1318 0 -1
Gyc2_1319 y2 0 x1319 0 1
Gyc2_1320 y2 0 x1320 0 1
Gyc2_1321 y2 0 x1321 0 -1
Gyc2_1322 y2 0 x1322 0 1
Gyc2_1323 y2 0 x1323 0 -1
Gyc2_1324 y2 0 x1324 0 1
Gyc2_1325 y2 0 x1325 0 -1
Gyc2_1326 y2 0 x1326 0 1
Gyc2_1327 y2 0 x1327 0 -1
Gyc2_1328 y2 0 x1328 0 -1
Gyc2_1329 y2 0 x1329 0 1
Gyc2_1330 y2 0 x1330 0 1
Gyc2_1331 y2 0 x1331 0 -1
Gyc2_1332 y2 0 x1332 0 -1
Gyc2_1333 y2 0 x1333 0 1
Gyc2_1334 y2 0 x1334 0 1
Gyc2_1335 y2 0 x1335 0 -1
Gyc2_1336 y2 0 x1336 0 -1
Gyc2_1337 y2 0 x1337 0 1
Gyc2_1338 y2 0 x1338 0 -1
Gyc2_1339 y2 0 x1339 0 1
Gyc2_1340 y2 0 x1340 0 1
Gyc2_1341 y2 0 x1341 0 1
Gyc2_1342 y2 0 x1342 0 -1
Gyc2_1343 y2 0 x1343 0 1
Gyc2_1344 y2 0 x1344 0 1
Gyc2_1345 y2 0 x1345 0 -1
Gyc2_1346 y2 0 x1346 0 -1
Gyc2_1347 y2 0 x1347 0 -1
Gyc2_1348 y2 0 x1348 0 -1
Gyc2_1349 y2 0 x1349 0 1
Gyc2_1350 y2 0 x1350 0 1
Gyc2_1351 y2 0 x1351 0 -1
Gyc2_1352 y2 0 x1352 0 1
Gyc2_1353 y2 0 x1353 0 -1
Gyc2_1354 y2 0 x1354 0 1
Gyc2_1355 y2 0 x1355 0 1
Gyc2_1356 y2 0 x1356 0 -1
Gyc2_1357 y2 0 x1357 0 -1
Gyc2_1358 y2 0 x1358 0 -1
Gyc2_1359 y2 0 x1359 0 1
Gyc2_1360 y2 0 x1360 0 -1
Gyc2_1361 y2 0 x1361 0 -1
Gyc2_1362 y2 0 x1362 0 1
Gyc2_1363 y2 0 x1363 0 -1
Gyc2_1364 y2 0 x1364 0 1
Gyc2_1365 y2 0 x1365 0 -1
Gyc2_1366 y2 0 x1366 0 -1
Gyc2_1367 y2 0 x1367 0 1
Gyc2_1368 y2 0 x1368 0 1
Gyc2_1369 y2 0 x1369 0 -1
Gyc2_1370 y2 0 x1370 0 -1
Gyc2_1371 y2 0 x1371 0 1
Gyc2_1372 y2 0 x1372 0 1
Gyc2_1373 y2 0 x1373 0 -1
Gyc2_1374 y2 0 x1374 0 -1
Gyc2_1375 y2 0 x1375 0 1
Gyc2_1376 y2 0 x1376 0 1
Gyc2_1377 y2 0 x1377 0 1
Gyc2_1378 y2 0 x1378 0 1
Gyc2_1379 y2 0 x1379 0 -1
Gyc2_1380 y2 0 x1380 0 -1
Gyc2_1381 y2 0 x1381 0 1
Gyc2_1382 y2 0 x1382 0 1
Gyc2_1383 y2 0 x1383 0 -1
Gyc2_1384 y2 0 x1384 0 -1
Gyc2_1385 y2 0 x1385 0 -1
Gyc2_1386 y2 0 x1386 0 1
Gyc2_1387 y2 0 x1387 0 -1
Gyc2_1388 y2 0 x1388 0 1
Gyc2_1389 y2 0 x1389 0 1
Gyc2_1390 y2 0 x1390 0 -1
Gyc2_1391 y2 0 x1391 0 -1
Gyc2_1392 y2 0 x1392 0 1
Gyc2_1393 y2 0 x1393 0 1
Gyc2_1394 y2 0 x1394 0 -1
Gyc2_1395 y2 0 x1395 0 -1
Gyc2_1396 y2 0 x1396 0 -1
Gyc2_1397 y2 0 x1397 0 -1
Gyc2_1398 y2 0 x1398 0 1
Gyc2_1399 y2 0 x1399 0 -1
Gyc2_1400 y2 0 x1400 0 1
Gyc2_1401 y2 0 x1401 0 -1
Gyc2_1402 y2 0 x1402 0 -1
Gyc2_1403 y2 0 x1403 0 -1
Gyc2_1404 y2 0 x1404 0 -1
Gyc2_1405 y2 0 x1405 0 1
Gyc2_1406 y2 0 x1406 0 1
Gyc2_1407 y2 0 x1407 0 -1
Gyc2_1408 y2 0 x1408 0 1
Gyc2_1409 y2 0 x1409 0 1
Gyc2_1410 y2 0 x1410 0 1
Gyc2_1411 y2 0 x1411 0 1
Gyc2_1412 y2 0 x1412 0 1
Gyc2_1413 y2 0 x1413 0 -1
Gyc2_1414 y2 0 x1414 0 -1
Gyc2_1415 y2 0 x1415 0 1
Gyc2_1416 y2 0 x1416 0 -1
Gyc2_1417 y2 0 x1417 0 -1
Gyc2_1418 y2 0 x1418 0 -1
Gyc2_1419 y2 0 x1419 0 1
Gyc2_1420 y2 0 x1420 0 -1
Gyc2_1421 y2 0 x1421 0 1
Gyc2_1422 y2 0 x1422 0 -1
Gyc2_1423 y2 0 x1423 0 1
Gyc2_1424 y2 0 x1424 0 1
Gyc2_1425 y2 0 x1425 0 -1
Gyc2_1426 y2 0 x1426 0 -1
Gyc2_1427 y2 0 x1427 0 -1
Gyc2_1428 y2 0 x1428 0 -1
Gyc2_1429 y2 0 x1429 0 1
Gyc2_1430 y2 0 x1430 0 1
Gyc2_1431 y2 0 x1431 0 1
Gyc2_1432 y2 0 x1432 0 1
Gyc2_1433 y2 0 x1433 0 -1
Gyc2_1434 y2 0 x1434 0 1
Gyc2_1435 y2 0 x1435 0 1
Gyc2_1436 y2 0 x1436 0 -1
Gyc2_1437 y2 0 x1437 0 -1
Gyc2_1438 y2 0 x1438 0 1
Gyc2_1439 y2 0 x1439 0 -1
Gyc2_1440 y2 0 x1440 0 -1
Gyc2_1441 y2 0 x1441 0 -1
Gyc2_1442 y2 0 x1442 0 -1
Gyc2_1443 y2 0 x1443 0 1
Gyc2_1444 y2 0 x1444 0 -1
Gyc2_1445 y2 0 x1445 0 1
Gyc2_1446 y2 0 x1446 0 -1
Gyc2_1447 y2 0 x1447 0 -1
Gyc2_1448 y2 0 x1448 0 -1
Gyc2_1449 y2 0 x1449 0 -1
Gyc2_1450 y2 0 x1450 0 1
Gyc2_1451 y2 0 x1451 0 -1
Gyc2_1452 y2 0 x1452 0 -1
Gyc2_1453 y2 0 x1453 0 -0.250929404461565
Gyc2_1454 y2 0 x1454 0 -1
Gyc2_1455 y2 0 x1455 0 -1
Gyc2_1456 y2 0 x1456 0 -1
Gyc2_1457 y2 0 x1457 0 1
Gyc2_1458 y2 0 x1458 0 -1
Gyc2_1459 y2 0 x1459 0 -1
Gyc2_1460 y2 0 x1460 0 1
Gyc2_1461 y2 0 x1461 0 1
Gyc2_1462 y2 0 x1462 0 -1
Gyc2_1463 y2 0 x1463 0 1
Gyc2_1464 y2 0 x1464 0 -1
Gyc2_1465 y2 0 x1465 0 -1
Gyc2_1466 y2 0 x1466 0 1
Gyc2_1467 y2 0 x1467 0 1
Gyc2_1468 y2 0 x1468 0 -1
Gyc2_1469 y2 0 x1469 0 1
Gyc2_1470 y2 0 x1470 0 -1
Gyc2_1471 y2 0 x1471 0 -1
Gyc2_1472 y2 0 x1472 0 -1
Gyc2_1473 y2 0 x1473 0 1
Gyc2_1474 y2 0 x1474 0 -1
Gyc2_1475 y2 0 x1475 0 -1
Gyc2_1476 y2 0 x1476 0 1
Gyc2_1477 y2 0 x1477 0 1
Gyc2_1478 y2 0 x1478 0 1
Gyc2_1479 y2 0 x1479 0 -1
Gyc2_1480 y2 0 x1480 0 1
Gyc2_1481 y2 0 x1481 0 -1
Gyc2_1482 y2 0 x1482 0 1
Gyc2_1483 y2 0 x1483 0 1
Gyc2_1484 y2 0 x1484 0 -1
Gyc2_1485 y2 0 x1485 0 1
Gyc2_1486 y2 0 x1486 0 1
Gyc2_1487 y2 0 x1487 0 1
Gyc2_1488 y2 0 x1488 0 1
Gyc2_1489 y2 0 x1489 0 -1
Gyc2_1490 y2 0 x1490 0 1
Gyc2_1491 y2 0 x1491 0 -1
Gyc2_1492 y2 0 x1492 0 1
Gyc2_1493 y2 0 x1493 0 -1
Gyc2_1494 y2 0 x1494 0 1
Gyc2_1495 y2 0 x1495 0 1
Gyc2_1496 y2 0 x1496 0 -1
Gyc2_1497 y2 0 x1497 0 1
Gyc2_1498 y2 0 x1498 0 -1
Gyc2_1499 y2 0 x1499 0 -1
Gyc2_1500 y2 0 x1500 0 -1
Gyc2_1501 y2 0 x1501 0 1
Gyc2_1502 y2 0 x1502 0 1
Gyc2_1503 y2 0 x1503 0 -1
Gyc2_1504 y2 0 x1504 0 -1
Gyc2_1505 y2 0 x1505 0 -1
Gyc2_1506 y2 0 x1506 0 -1
Gyc2_1507 y2 0 x1507 0 1
Gyc2_1508 y2 0 x1508 0 -1
Gyc2_1509 y2 0 x1509 0 1
Gyc2_1510 y2 0 x1510 0 -1
Gyc2_1511 y2 0 x1511 0 1
Gyc2_1512 y2 0 x1512 0 -1
Gyc2_1513 y2 0 x1513 0 -1
Gyc2_1514 y2 0 x1514 0 -1
Gyc2_1515 y2 0 x1515 0 1
Gyc2_1516 y2 0 x1516 0 -1
Gyc2_1517 y2 0 x1517 0 1
Gyc2_1518 y2 0 x1518 0 1
Gyc2_1519 y2 0 x1519 0 -1
Gyc2_1520 y2 0 x1520 0 -1
Gyc2_1521 y2 0 x1521 0 -1
Gyc2_1522 y2 0 x1522 0 1
Gyc2_1523 y2 0 x1523 0 1
Gyc2_1524 y2 0 x1524 0 -1
Gyc2_1525 y2 0 x1525 0 -1
Gyc2_1526 y2 0 x1526 0 -1
Gyc2_1527 y2 0 x1527 0 -1
Gyc2_1528 y2 0 x1528 0 1
Gyc2_1529 y2 0 x1529 0 -1
Gyc2_1530 y2 0 x1530 0 -1
Gyc2_1531 y2 0 x1531 0 1
Gyc2_1532 y2 0 x1532 0 -1
Gyc2_1533 y2 0 x1533 0 1
Gyc2_1534 y2 0 x1534 0 1
Gyc2_1535 y2 0 x1535 0 1
Gyc2_1536 y2 0 x1536 0 1
Gyc2_1537 y2 0 x1537 0 -1
Gyc2_1538 y2 0 x1538 0 1
Gyc2_1539 y2 0 x1539 0 1
Gyc2_1540 y2 0 x1540 0 1
Gyc2_1541 y2 0 x1541 0 1
Gyc2_1542 y2 0 x1542 0 1
Gyc2_1543 y2 0 x1543 0 -1
Gyc2_1544 y2 0 x1544 0 1
Gyc2_1545 y2 0 x1545 0 1
Gyc2_1546 y2 0 x1546 0 -1
Gyc2_1547 y2 0 x1547 0 -1
Gyc2_1548 y2 0 x1548 0 -1
Gyc2_1549 y2 0 x1549 0 -1
Gyc2_1550 y2 0 x1550 0 -1
Gyc2_1551 y2 0 x1551 0 -0.874267151697707
Gyc2_1552 y2 0 x1552 0 -1
Gyc2_1553 y2 0 x1553 0 -1
Gyc2_1554 y2 0 x1554 0 -1
Gyc2_1555 y2 0 x1555 0 1
Gyc2_1556 y2 0 x1556 0 1
Gyc2_1557 y2 0 x1557 0 -1
Gyc2_1558 y2 0 x1558 0 1
Gyc2_1559 y2 0 x1559 0 1
Gyc2_1560 y2 0 x1560 0 1
Gyc2_1561 y2 0 x1561 0 -1
Gyc2_1562 y2 0 x1562 0 1
Gyc2_1563 y2 0 x1563 0 -1
Gyc2_1564 y2 0 x1564 0 -1
Gyc2_1565 y2 0 x1565 0 -1
Gyc2_1566 y2 0 x1566 0 1
Gyc2_1567 y2 0 x1567 0 1
Gyc2_1568 y2 0 x1568 0 -1
Gyc2_1569 y2 0 x1569 0 1
Gyc2_1570 y2 0 x1570 0 1
Gyc2_1571 y2 0 x1571 0 -1
Gyc2_1572 y2 0 x1572 0 1
Gyc2_1573 y2 0 x1573 0 1
Gyc2_1574 y2 0 x1574 0 1
Gyc2_1575 y2 0 x1575 0 1
Gyc2_1576 y2 0 x1576 0 1
Gyc2_1577 y2 0 x1577 0 1
Gyc2_1578 y2 0 x1578 0 -1
Gyc2_1579 y2 0 x1579 0 1
Gyc2_1580 y2 0 x1580 0 1
Gyc2_1581 y2 0 x1581 0 -1
Gyc2_1582 y2 0 x1582 0 1
Gyc2_1583 y2 0 x1583 0 1
Gyc2_1584 y2 0 x1584 0 1
Gyc2_1585 y2 0 x1585 0 -1
Gyc2_1586 y2 0 x1586 0 1
Gyc2_1587 y2 0 x1587 0 -1
Gyc2_1588 y2 0 x1588 0 -1
Gyc2_1589 y2 0 x1589 0 -1
Gyc2_1590 y2 0 x1590 0 -1
Gyc2_1591 y2 0 x1591 0 -1
Gyc2_1592 y2 0 x1592 0 -1
Gyc2_1593 y2 0 x1593 0 -1
Gyc2_1594 y2 0 x1594 0 -1
Gyc2_1595 y2 0 x1595 0 1
Gyc2_1596 y2 0 x1596 0 -1
Gyc2_1597 y2 0 x1597 0 -1
Gyc2_1598 y2 0 x1598 0 1
Gyc2_1599 y2 0 x1599 0 1
Gyc2_1600 y2 0 x1600 0 -1
Gyc2_1601 y2 0 x1601 0 1
Gyc2_1602 y2 0 x1602 0 -1
.ENDS
