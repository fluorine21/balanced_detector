* Equivalent circuit model for CMA-5043+_5V_Plus25DegC.ckt
.SUBCKT CMA-5043+_5V_Plus25DegC po1 po2
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Vsp2 po2 p2 0
Vsr2 p2 pr2 0
Rp2 pr2 0 50
Ru2 u2 0 50
Fr2 u2 0 Vsr2 -1
Fu2 u2 0 Vsp2 -1
Ry2 y2 0 1
Gy2 p2 0 y2 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 2.09429757386434
Cx1 x1 xm1 2.87060508922215e-13
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.000149951069880376
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -445.251537372569
Cx2 x2 xm2 2.87060508922216e-13
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.0667659443948988
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 37.7178314529486
Cx3 x3 xm3 2.14951724198048e-13
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -0.000104470432497296
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -48.8139755625609
Cx4 x4 xm4 2.14951724198048e-13
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 0.00509961713893317
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 3.90299552268256
Cx5 x5 xm5 2.64800814690544e-13
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -2.23795403791762e-05
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -335.499699936289
Cx6 x6 xm6 2.64800814690544e-13
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 0.00750832908192567
Rx7 x7 0 1
Fxc7_8 x7 0 Vx8 24.6178887893632
Cx7 x7 xm7 9.06783631436284e-13
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 -0.0283470144271603
Rx8 x8 0 1
Fxc8_7 x8 0 Vx7 -4.99671192362294
Cx8 x8 xm8 9.06783631436284e-13
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 0.141641864987303
Rx9 x9 0 1
Fxc9_10 x9 0 Vx10 28.8495040748833
Cx9 x9 xm9 3.37827865050702e-13
Vx9 xm9 0 0
Gx9_1 x9 0 u1 0 -0.000457376606440122
Rx10 x10 0 1
Fxc10_9 x10 0 Vx9 -33.4199174509494
Cx10 x10 xm10 3.37827865050702e-13
Vx10 xm10 0 0
Gx10_1 x10 0 u1 0 0.0152854884312242
Rx11 x11 0 1
Fxc11_12 x11 0 Vx12 36.3267548797069
Cx11 x11 xm11 2.16746118370639e-13
Vx11 xm11 0 0
Gx11_1 x11 0 u1 0 -0.000119108042850154
Rx12 x12 0 1
Fxc12_11 x12 0 Vx11 -67.0292088175732
Cx12 x12 xm12 2.16746118370639e-13
Vx12 xm12 0 0
Gx12_1 x12 0 u1 0 0.00798371787605541
Rx13 x13 0 1
Fxc13_14 x13 0 Vx14 52.0091341880116
Cx13 x13 xm13 2.35673728092649e-13
Vx13 xm13 0 0
Gx13_1 x13 0 u1 0 -2.78539292500512e-05
Rx14 x14 0 1
Fxc14_13 x14 0 Vx13 -44.3284359836786
Cx14 x14 xm14 2.35673728092649e-13
Vx14 xm14 0 0
Gx14_1 x14 0 u1 0 0.00123472111965481
Rx15 x15 0 1
Fxc15_16 x15 0 Vx16 9.61549107737617
Cx15 x15 xm15 9.9938565516691e-13
Vx15 xm15 0 0
Gx15_1 x15 0 u1 0 -0.0132320427207703
Rx16 x16 0 1
Fxc16_15 x16 0 Vx15 -14.2569754549145
Cx16 x16 xm16 9.9938565516691e-13
Vx16 xm16 0 0
Gx16_1 x16 0 u1 0 0.188648908288402
Rx17 x17 0 1
Fxc17_18 x17 0 Vx18 27.2894618266908
Cx17 x17 xm17 1.58482941113653e-13
Vx17 xm17 0 0
Gx17_1 x17 0 u1 0 -4.33500658190099e-06
Rx18 x18 0 1
Fxc18_17 x18 0 Vx17 -222.530142256075
Cx18 x18 xm18 1.58482941113653e-13
Vx18 xm18 0 0
Gx18_1 x18 0 u1 0 0.000964669631351448
Rx19 x19 0 1
Fxc19_20 x19 0 Vx20 15.509033142785
Cx19 x19 xm19 2.96947443018644e-13
Vx19 xm19 0 0
Gx19_1 x19 0 u1 0 -3.37955711355307e-05
Rx20 x20 0 1
Fxc20_19 x20 0 Vx19 -116.04935477903
Cx20 x20 xm20 2.96947443018644e-13
Vx20 xm20 0 0
Gx20_1 x20 0 u1 0 0.00392195422466717
Rx21 x21 0 1
Fxc21_22 x21 0 Vx22 46.5001671964016
Cx21 x21 xm21 2.82489214445738e-13
Vx21 xm21 0 0
Gx21_1 x21 0 u1 0 -2.0017229602428e-05
Rx22 x22 0 1
Fxc22_21 x22 0 Vx21 -47.8089659008142
Cx22 x22 xm22 2.82489214445738e-13
Vx22 xm22 0 0
Gx22_1 x22 0 u1 0 0.00095700304749125
Rx23 x23 0 1
Fxc23_24 x23 0 Vx24 29.3265475148589
Cx23 x23 xm23 1.25157800297801e-12
Vx23 xm23 0 0
Gx23_1 x23 0 u1 0 -0.0103140208552761
Rx24 x24 0 1
Fxc24_23 x24 0 Vx23 -4.22305594485865
Cx24 x24 xm24 1.25157800297801e-12
Vx24 xm24 0 0
Gx24_1 x24 0 u1 0 0.04355668708827
Rx25 x25 0 1
Fxc25_26 x25 0 Vx26 21.7082997240386
Cx25 x25 xm25 1.51094605540703e-12
Vx25 xm25 0 0
Gx25_1 x25 0 u1 0 -0.0115929926047637
Rx26 x26 0 1
Fxc26_25 x26 0 Vx25 -4.58115378939401
Cx26 x26 xm26 1.51094605540703e-12
Vx26 xm26 0 0
Gx26_1 x26 0 u1 0 0.0531092820017299
Rx27 x27 0 1
Fxc27_28 x27 0 Vx28 1.40522799907503
Cx27 x27 xm27 1.70972884859627e-12
Vx27 xm27 0 0
Gx27_1 x27 0 u1 0 -0.000772671018570193
Rx28 x28 0 1
Fxc28_27 x28 0 Vx27 -64.4081824157388
Cx28 x28 xm28 1.70972884859627e-12
Vx28 xm28 0 0
Gx28_1 x28 0 u1 0 0.0497663359114237
Rx29 x29 0 1
Fxc29_30 x29 0 Vx30 0.624885741261362
Cx29 x29 xm29 1.61515298397391e-12
Vx29 xm29 0 0
Gx29_1 x29 0 u1 0 -0.000256334467977839
Rx30 x30 0 1
Fxc30_29 x30 0 Vx29 -250.070669835055
Cx30 x30 xm30 1.61515298397391e-12
Vx30 xm30 0 0
Gx30_1 x30 0 u1 0 0.0641017321090306
Rx31 x31 0 1
Fxc31_32 x31 0 Vx32 1.72945456140906
Cx31 x31 xm31 3.3832600882424e-12
Vx31 xm31 0 0
Gx31_1 x31 0 u1 0 -0.0121248297230833
Rx32 x32 0 1
Fxc32_31 x32 0 Vx31 -20.1948098501078
Cx32 x32 xm32 3.3832600882424e-12
Vx32 xm32 0 0
Gx32_1 x32 0 u1 0 0.244858630722602
Rx33 x33 0 1
Fxc33_34 x33 0 Vx34 12.2736156153286
Cx33 x33 xm33 6.36249392361281e-12
Vx33 xm33 0 0
Gx33_1 x33 0 u1 0 -0.146340705650046
Rx34 x34 0 1
Fxc34_33 x34 0 Vx33 -1.38675608761447
Cx34 x34 xm34 6.36249392361281e-12
Vx34 xm34 0 0
Gx34_1 x34 0 u1 0 0.202938864425998
Rx35 x35 0 1
Fxc35_36 x35 0 Vx36 7.25559809336935
Cx35 x35 xm35 4.08890323417608e-12
Vx35 xm35 0 0
Gx35_1 x35 0 u1 0 -0.00610556124133608
Rx36 x36 0 1
Fxc36_35 x36 0 Vx35 -7.33457076772417
Cx36 x36 xm36 4.08890323417608e-12
Vx36 xm36 0 0
Gx36_1 x36 0 u1 0 0.0447816710012533
Rx37 x37 0 1
Fxc37_38 x37 0 Vx38 22.5908294986345
Cx37 x37 xm37 1.41898003518717e-11
Vx37 xm37 0 0
Gx37_1 x37 0 u1 0 -0.234512886573611
Rx38 x38 0 1
Fxc38_37 x38 0 Vx37 -0.295661942189029
Cx38 x38 xm38 1.41898003518717e-11
Vx38 xm38 0 0
Gx38_1 x38 0 u1 0 0.0693365355127092
Rx39 x39 0 1
Fxc39_40 x39 0 Vx40 3.36171152527201
Cx39 x39 xm39 3.02223658791127e-11
Vx39 xm39 0 0
Gx39_1 x39 0 u1 0 -0.612257190887511
Rx40 x40 0 1
Fxc40_39 x40 0 Vx39 -0.73155948098281
Cx40 x40 xm40 3.02223658791127e-11
Vx40 xm40 0 0
Gx40_1 x40 0 u1 0 0.447902552793661
Rx41 x41 0 1
Fxc41_42 x41 0 Vx42 10.7468518171504
Cx41 x41 xm41 1.30273315544064e-11
Vx41 xm41 0 0
Gx41_1 x41 0 u1 0 -0.00425896546207179
Rx42 x42 0 1
Fxc42_41 x42 0 Vx41 -2.77463905341064
Cx42 x42 xm42 1.30273315544064e-11
Vx42 xm42 0 0
Gx42_1 x42 0 u1 0 0.0118170918981915
Rx43 x43 0 1
Fxc43_44 x43 0 Vx44 3.36434889032178
Cx43 x43 xm43 4.87133831260231e-12
Vx43 xm43 0 0
Gx43_1 x43 0 u1 0 -3.0121413672702e-05
Rx44 x44 0 1
Fxc44_43 x44 0 Vx43 -81.1455606399185
Cx44 x44 xm44 4.87133831260231e-12
Vx44 xm44 0 0
Gx44_1 x44 0 u1 0 0.00244421899973831
Rx45 x45 0 1
Fxc45_46 x45 0 Vx46 1.61998700601747
Cx45 x45 xm45 7.06557064659634e-11
Vx45 xm45 0 0
Gx45_1 x45 0 u1 0 -0.744361500392355
Rx46 x46 0 1
Fxc46_45 x46 0 Vx45 -0.932110779964664
Cx46 x46 xm46 7.06557064659634e-11
Vx46 xm46 0 0
Gx46_1 x46 0 u1 0 0.693827378706385
Rx47 x47 0 1
Fxc47_48 x47 0 Vx48 3.0556073611081
Cx47 x47 xm47 9.00586691578378e-12
Vx47 xm47 0 0
Gx47_1 x47 0 u1 0 -2.27633167309635e-05
Rx48 x48 0 1
Fxc48_47 x48 0 Vx47 -111.996144516901
Cx48 x48 xm48 9.00586691578377e-12
Vx48 xm48 0 0
Gx48_1 x48 0 u1 0 0.00254940371028497
Rx49 x49 0 1
Fxc49_50 x49 0 Vx50 209.066355813791
Cx49 x49 xm49 6.72924348226814e-13
Vx49 xm49 0 0
Gx49_1 x49 0 u1 0 -1.72848174119649e-07
Rx50 x50 0 1
Fxc50_49 x50 0 Vx49 -303.5846766105
Cx50 x50 xm50 6.72924348226814e-13
Vx50 xm50 0 0
Gx50_1 x50 0 u1 0 5.24740570428291e-05
Rx51 x51 0 1
Fxc51_52 x51 0 Vx52 14.2532269714476
Cx51 x51 xm51 7.40586010206479e-13
Vx51 xm51 0 0
Gx51_1 x51 0 u1 0 -1.63982640887449e-08
Rx52 x52 0 1
Fxc52_51 x52 0 Vx51 -4179.62689532179
Cx52 x52 xm52 7.40586010206479e-13
Vx52 xm52 0 0
Gx52_1 x52 0 u1 0 6.85386256219076e-05
Rx53 x53 0 1
Fxc53_54 x53 0 Vx54 0.0534208873918435
Cx53 x53 xm53 2.7189670410967e-10
Vx53 xm53 0 0
Gx53_1 x53 0 u1 0 -16.7327745838584
Rx54 x54 0 1
Fxc54_53 x54 0 Vx53 -0.11560606544592
Cx54 x54 xm54 2.7189670410967e-10
Vx54 xm54 0 0
Gx54_1 x54 0 u1 0 1.93441023363336
Rx55 x55 0 1
Fxc55_56 x55 0 Vx56 75.6700575339533
Cx55 x55 xm55 3.40336796714079e-13
Vx55 xm55 0 0
Gx55_1 x55 0 u1 0 -1.14949252259274e-08
Rx56 x56 0 1
Fxc56_55 x56 0 Vx55 -4273.80783317262
Cx56 x56 xm56 3.40336796714079e-13
Vx56 xm56 0 0
Gx56_1 x56 0 u1 0 4.91271014723022e-05
Rx57 x57 0 1
Fxc57_58 x57 0 Vx58 7.91486403926958
Cx57 x57 xm57 1.77838009044698e-11
Vx57 xm57 0 0
Gx57_1 x57 0 u1 0 -0.000599939984699646
Rx58 x58 0 1
Fxc58_57 x58 0 Vx57 -16.0224274862753
Cx58 x58 xm58 1.77838009044698e-11
Vx58 xm58 0 0
Gx58_1 x58 0 u1 0 0.00961249490096718
Rx59 x59 0 1
Fxc59_60 x59 0 Vx60 6607.97178609309
Cx59 x59 xm59 6.45459166206642e-14
Vx59 xm59 0 0
Gx59_1 x59 0 u1 0 -6.45789721874064e-09
Rx60 x60 0 1
Fxc60_59 x60 0 Vx59 -1519.52832514805
Cx60 x60 xm60 6.45459166206642e-14
Vx60 xm60 0 0
Gx60_1 x60 0 u1 0 9.81295774477122e-06
Rx61 x61 0 1
Fxc61_62 x61 0 Vx62 31.3672180629436
Cx61 x61 xm61 3.60587813907164e-12
Vx61 xm61 0 0
Gx61_1 x61 0 u1 0 -7.06813193854952e-06
Rx62 x62 0 1
Fxc62_61 x62 0 Vx61 -108.198098019568
Cx62 x62 xm62 3.60587813907164e-12
Vx62 xm62 0 0
Gx62_1 x62 0 u1 0 0.000764758432302417
Rx63 x63 0 1
Fxc63_64 x63 0 Vx64 0.970794556404795
Cx63 x63 xm63 1.33799391561211e-11
Vx63 xm63 0 0
Gx63_1 x63 0 u1 0 -7.02762529848386e-05
Rx64 x64 0 1
Fxc64_63 x64 0 Vx63 -293.307078040876
Cx64 x64 xm64 1.33799391561211e-11
Vx64 xm64 0 0
Gx64_1 x64 0 u1 0 0.0206125224186444
Rx65 x65 0 1
Fxc65_66 x65 0 Vx66 140.74212076884
Cx65 x65 xm65 2.86431819527606e-12
Vx65 xm65 0 0
Gx65_1 x65 0 u1 0 -8.29427267619837e-06
Rx66 x66 0 1
Fxc66_65 x66 0 Vx65 -41.0983957834867
Cx66 x66 xm66 2.86431819527606e-12
Vx66 xm66 0 0
Gx66_1 x66 0 u1 0 0.00034088130118256
Rx67 x67 0 1
Fxc67_68 x67 0 Vx68 101.574703323604
Cx67 x67 xm67 7.0808537117008e-12
Vx67 xm67 0 0
Gx67_1 x67 0 u1 0 -0.000134357302801061
Rx68 x68 0 1
Fxc68_67 x68 0 Vx67 -10.6013913438328
Cx68 x68 xm68 7.0808537117008e-12
Vx68 xm68 0 0
Gx68_1 x68 0 u1 0 0.00142437434689589
Rx69 x69 0 1
Fxc69_70 x69 0 Vx70 32.5244512511448
Cx69 x69 xm69 8.39484573603046e-12
Vx69 xm69 0 0
Gx69_1 x69 0 u1 0 -6.16257352745165e-05
Rx70 x70 0 1
Fxc70_69 x70 0 Vx69 -26.5921344226316
Cx70 x70 xm70 8.39484573603046e-12
Vx70 xm70 0 0
Gx70_1 x70 0 u1 0 0.00163875983631345
Rx71 x71 0 1
Fxc71_72 x71 0 Vx72 1597.17633201235
Cx71 x71 xm71 2.83045279415423e-13
Vx71 xm71 0 0
Gx71_1 x71 0 u1 0 -7.78590865211595e-08
Rx72 x72 0 1
Fxc72_71 x72 0 Vx71 -501.488167164467
Cx72 x72 xm72 2.83045279415423e-13
Vx72 xm72 0 0
Gx72_1 x72 0 u1 0 3.9045410596596e-05
Rx73 x73 0 1
Fxc73_74 x73 0 Vx74 163.081677433848
Cx73 x73 xm73 5.19274272676225e-12
Vx73 xm73 0 0
Gx73_1 x73 0 u1 0 -1.2410753407805e-05
Rx74 x74 0 1
Fxc74_73 x74 0 Vx73 -16.5231311120809
Cx74 x74 xm74 5.19274272676225e-12
Vx74 xm74 0 0
Gx74_1 x74 0 u1 0 0.000205064505756866
Rx75 x75 0 1
Fxc75_76 x75 0 Vx76 562.687535923902
Cx75 x75 xm75 6.76962091359381e-13
Vx75 xm75 0 0
Gx75_1 x75 0 u1 0 -9.29785289638722e-08
Rx76 x76 0 1
Fxc76_75 x76 0 Vx75 -305.328657198455
Cx76 x76 xm76 6.76962091359381e-13
Vx76 xm76 0 0
Gx76_1 x76 0 u1 0 2.83890093968268e-05
Rx77 x77 0 1
Fxc77_78 x77 0 Vx78 110.355496324475
Cx77 x77 xm77 1.60390660485385e-11
Vx77 xm77 0 0
Gx77_1 x77 0 u1 0 -0.000251629984138903
Rx78 x78 0 1
Fxc78_77 x78 0 Vx77 -2.85603597824502
Cx78 x78 xm78 1.60390660485385e-11
Vx78 xm78 0 0
Gx78_1 x78 0 u1 0 0.00071866428790593
Rx79 x79 0 1
Fxc79_80 x79 0 Vx80 0.524658073787078
Cx79 x79 xm79 3.65373015413682e-11
Vx79 xm79 0 0
Gx79_1 x79 0 u1 0 -0.000209006807996916
Rx80 x80 0 1
Fxc80_79 x80 0 Vx79 -131.971525733187
Cx80 x80 xm80 3.65373015413682e-11
Vx80 xm80 0 0
Gx80_1 x80 0 u1 0 0.0275829473399762
Rx81 x81 0 1
Fxc81_82 x81 0 Vx82 98.3615319636901
Cx81 x81 xm81 4.9605444448296e-12
Vx81 xm81 0 0
Gx81_1 x81 0 u1 0 -4.79488153908484e-06
Rx82 x82 0 1
Fxc82_81 x82 0 Vx81 -46.7618718670489
Cx82 x82 xm82 4.9605444448296e-12
Vx82 xm82 0 0
Gx82_1 x82 0 u1 0 0.000224217636148364
Rx83 x83 0 1
Fxc83_84 x83 0 Vx84 20.0398020738261
Cx83 x83 xm83 1.85213203877505e-12
Vx83 xm83 0 0
Gx83_1 x83 0 u1 0 -1.19023975072567e-07
Rx84 x84 0 1
Fxc84_83 x84 0 Vx83 -1836.7047721807
Cx84 x84 xm84 1.85213203877505e-12
Vx84 xm84 0 0
Gx84_1 x84 0 u1 0 0.000218611903019701
Rx85 x85 0 1
Fxc85_86 x85 0 Vx86 44.6077650092189
Cx85 x85 xm85 6.12244434678794e-12
Vx85 xm85 0 0
Gx85_1 x85 0 u1 0 -4.96508506633859e-06
Rx86 x86 0 1
Fxc86_85 x86 0 Vx85 -88.2816856942824
Cx86 x86 xm86 6.12244434678794e-12
Vx86 xm86 0 0
Gx86_1 x86 0 u1 0 0.000438326079271879
Rx87 x87 0 1
Fxc87_88 x87 0 Vx88 1181.89300944629
Cx87 x87 xm87 1.14029529690273e-12
Vx87 xm87 0 0
Gx87_1 x87 0 u1 0 -2.72230189976552e-07
Rx88 x88 0 1
Fxc88_87 x88 0 Vx87 -110.858410576864
Cx88 x88 xm88 1.14029529690273e-12
Vx88 xm88 0 0
Gx88_1 x88 0 u1 0 3.01790061718382e-05
Rx89 x89 0 1
Fxc89_90 x89 0 Vx90 491.969098447874
Cx89 x89 xm89 9.47069571391727e-12
Vx89 xm89 0 0
Gx89_1 x89 0 u1 0 -2.32713353055471e-05
Rx90 x90 0 1
Fxc90_89 x90 0 Vx89 -4.29840114567481
Cx90 x90 xm90 9.47069571391727e-12
Vx90 xm90 0 0
Gx90_1 x90 0 u1 0 0.000100029534338746
Rx91 x91 0 1
Fxc91_92 x91 0 Vx92 669.96282077103
Cx91 x91 xm91 1.41828331495617e-12
Vx91 xm91 0 0
Gx91_1 x91 0 u1 0 -7.30697663613735e-07
Rx92 x92 0 1
Fxc92_91 x92 0 Vx91 -151.199218134516
Cx92 x92 xm92 1.41828331495617e-12
Vx92 xm92 0 0
Gx92_1 x92 0 u1 0 0.000110480915431114
Rx93 x93 0 1
Fxc93_94 x93 0 Vx94 19.1597939071029
Cx93 x93 xm93 5.0878616870562e-12
Vx93 xm93 0 0
Gx93_1 x93 0 u1 0 -1.2518653813256e-06
Rx94 x94 0 1
Fxc94_93 x94 0 Vx93 -495.963972077337
Cx94 x94 xm94 5.0878616870562e-12
Vx94 xm94 0 0
Gx94_1 x94 0 u1 0 0.000620880127028355
Rx95 x95 0 1
Fxc95_96 x95 0 Vx96 7.86886673399765
Cx95 x95 xm95 4.66368852903178e-11
Vx95 xm95 0 0
Gx95_1 x95 0 u1 0 -0.000416736740754939
Rx96 x96 0 1
Fxc96_95 x96 0 Vx95 -18.5487607854936
Cx96 x96 xm96 4.66368852903178e-11
Vx96 xm96 0 0
Gx96_1 x96 0 u1 0 0.00772995011478962
Rx97 x97 0 1
Fxc97_98 x97 0 Vx98 46.57273051496
Cx97 x97 xm97 5.38073810888037e-12
Vx97 xm97 0 0
Gx97_1 x97 0 u1 0 -2.31248695644155e-06
Rx98 x98 0 1
Fxc98_97 x98 0 Vx97 -209.916194643155
Cx98 x98 xm98 5.38073810888037e-12
Vx98 xm98 0 0
Gx98_1 x98 0 u1 0 0.000485428462058141
Rx99 x99 0 1
Fxc99_100 x99 0 Vx100 154.621180355707
Cx99 x99 xm99 9.45572193374133e-12
Vx99 xm99 0 0
Gx99_1 x99 0 u1 0 -1.1762885680728e-05
Rx100 x100 0 1
Fxc100_99 x100 0 Vx99 -25.9316030607337
Cx100 x100 xm100 9.45572193374133e-12
Vx100 xm100 0 0
Gx100_1 x100 0 u1 0 0.000305030482321426
Rx101 x101 0 1
Fxc101_102 x101 0 Vx102 67.267513755542
Cx101 x101 xm101 1.20602139754355e-11
Vx101 xm101 0 0
Gx101_1 x101 0 u1 0 -1.69572574954266e-05
Rx102 x102 0 1
Fxc102_101 x102 0 Vx101 -43.9565752106921
Cx102 x102 xm102 1.20602139754355e-11
Vx102 xm102 0 0
Gx102_1 x102 0 u1 0 0.000745382964464792
Rx103 x103 0 1
Fxc103_104 x103 0 Vx104 244.134555454128
Cx103 x103 xm103 1.25498339510922e-11
Vx103 xm103 0 0
Gx103_1 x103 0 u1 0 -7.3931405139448e-06
Rx104 x104 0 1
Fxc104_103 x104 0 Vx103 -15.4411290431327
Cx104 x104 xm104 1.25498339510922e-11
Vx104 xm104 0 0
Gx104_1 x104 0 u1 0 0.000114158436709834
Rx105 x105 0 1
Fxc105_106 x105 0 Vx106 41.1219781367017
Cx105 x105 xm105 3.32631261202093e-11
Vx105 xm105 0 0
Gx105_1 x105 0 u1 0 -4.81356513856811e-05
Rx106 x106 0 1
Fxc106_105 x106 0 Vx105 -23.0543599215606
Cx106 x106 xm106 3.32631261202093e-11
Vx106 xm106 0 0
Gx106_1 x106 0 u1 0 0.00110973663210426
Rx107 x107 0 1
Fxc107_108 x107 0 Vx108 17.6320047809159
Cx107 x107 xm107 1.45379770932265e-10
Vx107 xm107 0 0
Gx107_1 x107 0 u1 0 -0.00137246973710192
Rx108 x108 0 1
Fxc108_107 x108 0 Vx107 -3.71520540693266
Cx108 x108 xm108 1.45379770932265e-10
Vx108 xm108 0 0
Gx108_1 x108 0 u1 0 0.00509900698813251
Rx109 x109 0 1
Fxc109_110 x109 0 Vx110 663.964978093968
Cx109 x109 xm109 4.64722716786655e-11
Vx109 xm109 0 0
Gx109_1 x109 0 u1 0 -6.16726235522221e-05
Rx110 x110 0 1
Fxc110_109 x110 0 Vx109 -4.942311054366
Cx110 x110 xm110 4.64722716786655e-11
Vx110 xm110 0 0
Gx110_1 x110 0 u1 0 0.0003048052891339
Rx111 x111 0 1
Fxc111_112 x111 0 Vx112 7.88054298013019
Cx111 x111 xm111 2.59641851055736e-10
Vx111 xm111 0 0
Gx111_1 x111 0 u1 0 -0.00039622983752322
Rx112 x112 0 1
Fxc112_111 x112 0 Vx111 -60.2028015819753
Cx112 x112 xm112 2.59641851055736e-10
Vx112 xm112 0 0
Gx112_1 x112 0 u1 0 0.0238541462892687
Rx113 x113 0 1
Fxc113_114 x113 0 Vx114 0.852015386400014
Cx113 x113 xm113 6.69011915274045e-09
Vx113 xm113 0 0
Gx113_1 x113 0 u1 0 -0.57375549423012
Rx114 x114 0 1
Fxc114_113 x114 0 Vx113 -5.85588652099324
Cx114 x114 xm114 6.69011915274045e-09
Vx114 xm114 0 0
Gx114_1 x114 0 u1 0 3.35984706500797
Rx115 x115 0 1
Fxc115_116 x115 0 Vx116 0.430281144205534
Cx115 x115 xm115 1.52744488718003e-09
Vx115 xm115 0 0
Gx115_1 x115 0 u1 0 -0.00464367320775955
Rx116 x116 0 1
Fxc116_115 x116 0 Vx115 -68.3212881669161
Cx116 x116 xm116 1.52744488718003e-09
Vx116 xm116 0 0
Gx116_1 x116 0 u1 0 0.317261735380328
Rx117 x117 0 1
Fxc117_118 x117 0 Vx118 41.6691319318108
Cx117 x117 xm117 1.70618985523348e-11
Vx117 xm117 0 0
Gx117_1 x117 0 u1 0 -4.87695569596373e-06
Rx118 x118 0 1
Fxc118_117 x118 0 Vx117 -836.822888292659
Cx118 x118 xm118 1.70618985523348e-11
Vx118 xm118 0 0
Gx118_1 x118 0 u1 0 0.0040811481515717
Rx119 x119 0 1
Cx119 x119 0 1.12913277439532e-08
Gx119_1 x119 0 u1 0 -0.960973157685528
Rx120 x120 0 1
Cx120 x120 0 2.13606987450335e-08
Gx120_1 x120 0 u1 0 -23.4069055687076
Rx121 x121 0 1
Fxc121_122 x121 0 Vx122 17.1392888247413
Cx121 x121 xm121 2.87060508922215e-13
Vx121 xm121 0 0
Gx121_2 x121 0 u2 0 -0.00111804352731375
Rx122 x122 0 1
Fxc122_121 x122 0 Vx121 -54.4065289997709
Cx122 x122 xm122 2.87060508922215e-13
Vx122 xm122 0 0
Gx122_2 x122 0 u2 0 0.0608288675918018
Rx123 x123 0 1
Fxc123_124 x123 0 Vx124 15.8654482460275
Cx123 x123 xm123 2.14951724198048e-13
Vx123 xm123 0 0
Gx123_2 x123 0 u2 0 -0.000153097712008718
Rx124 x124 0 1
Fxc124_123 x124 0 Vx123 -116.048237293139
Cx124 x124 xm124 2.14951724198049e-13
Vx124 xm124 0 0
Gx124_2 x124 0 u2 0 0.0177667196122244
Rx125 x125 0 1
Fxc125_126 x125 0 Vx126 180.861346752981
Cx125 x125 xm125 2.64800814690544e-13
Vx125 xm125 0 0
Gx125_2 x125 0 u2 0 -0.000656470906410051
Rx126 x126 0 1
Fxc126_125 x126 0 Vx125 -7.24009773354787
Cx126 x126 xm126 2.64800814690544e-13
Vx126 xm126 0 0
Gx126_2 x126 0 u2 0 0.00475291352163953
Rx127 x127 0 1
Fxc127_128 x127 0 Vx128 4.45923773022542
Cx127 x127 xm127 9.06783631436284e-13
Vx127 xm127 0 0
Gx127_2 x127 0 u2 0 -0.0069458033565874
Rx128 x128 0 1
Fxc128_127 x128 0 Vx127 -27.5850954557689
Cx128 x128 xm128 9.06783631436284e-13
Vx128 xm128 0 0
Gx128_2 x128 0 u2 0 0.191600648608463
Rx129 x129 0 1
Fxc129_130 x129 0 Vx130 74.5659867283274
Cx129 x129 xm129 3.37827865050702e-13
Vx129 xm129 0 0
Gx129_2 x129 0 u2 0 -0.00158120505896976
Rx130 x130 0 1
Fxc130_129 x130 0 Vx129 -12.9301319138469
Cx130 x130 xm130 3.37827865050702e-13
Vx130 xm130 0 0
Gx130_2 x130 0 u2 0 0.020445189995321
Rx131 x131 0 1
Fxc131_132 x131 0 Vx132 18.9430953366298
Cx131 x131 xm131 2.16746118370639e-13
Vx131 xm131 0 0
Gx131_2 x131 0 u2 0 -9.17545170976491e-05
Rx132 x132 0 1
Fxc132_131 x132 0 Vx131 -128.540430971081
Cx132 x132 xm132 2.16746118370639e-13
Vx132 xm132 0 0
Gx132_2 x132 0 u2 0 0.0117941651712753
Rx133 x133 0 1
Fxc133_134 x133 0 Vx134 19.2074583928036
Cx133 x133 xm133 2.35673728092649e-13
Vx133 xm133 0 0
Gx133_2 x133 0 u2 0 -3.54690720760159e-05
Rx134 x134 0 1
Fxc134_133 x134 0 Vx133 -120.030642694694
Cx134 x134 xm134 2.35673728092649e-13
Vx134 xm134 0 0
Gx134_2 x134 0 u2 0 0.00425737551706863
Rx135 x135 0 1
Fxc135_136 x135 0 Vx136 2.46192291029929
Cx135 x135 xm135 9.9938565516691e-13
Vx135 xm135 0 0
Gx135_2 x135 0 u2 0 -0.00404042205876885
Rx136 x136 0 1
Fxc136_135 x136 0 Vx135 -55.6832302520944
Cx136 x136 xm136 9.9938565516691e-13
Vx136 xm136 0 0
Gx136_2 x136 0 u2 0 0.224983751814067
Rx137 x137 0 1
Fxc137_138 x137 0 Vx138 231.557503081381
Cx137 x137 xm137 1.58482941113653e-13
Vx137 xm137 0 0
Gx137_2 x137 0 u2 0 -1.56541465454897e-05
Rx138 x138 0 1
Fxc138_137 x138 0 Vx137 -26.2255713659641
Cx138 x138 xm138 1.58482941113653e-13
Vx138 xm138 0 0
Gx138_2 x138 0 u2 0 0.000410538937402002
Rx139 x139 0 1
Fxc139_140 x139 0 Vx140 73.336272069362
Cx139 x139 xm139 2.96947443018644e-13
Vx139 xm139 0 0
Gx139_2 x139 0 u2 0 -0.00019608608592899
Rx140 x140 0 1
Fxc140_139 x140 0 Vx139 -24.5419250076487
Cx140 x140 xm140 2.96947443018644e-13
Vx140 xm140 0 0
Gx140_2 x140 0 u2 0 0.00481233001591264
Rx141 x141 0 1
Fxc141_142 x141 0 Vx142 25.8967253217752
Cx141 x141 xm141 2.82489214445738e-13
Vx141 xm141 0 0
Gx141_2 x141 0 u2 0 -1.7880123406017e-05
Rx142 x142 0 1
Fxc142_141 x142 0 Vx141 -85.8457924796235
Cx142 x142 xm142 2.82489214445738e-13
Vx142 xm142 0 0
Gx142_2 x142 0 u2 0 0.001534933363423
Rx143 x143 0 1
Fxc143_144 x143 0 Vx144 5.90482240736867
Cx143 x143 xm143 1.25157800297801e-12
Vx143 xm143 0 0
Gx143_2 x143 0 u2 0 -0.021421452301847
Rx144 x144 0 1
Fxc144_143 x144 0 Vx143 -20.9739840219842
Cx144 x144 xm144 1.25157800297801e-12
Vx144 xm144 0 0
Gx144_2 x144 0 u2 0 0.449293198306636
Rx145 x145 0 1
Fxc145_146 x145 0 Vx146 75.1311877867193
Cx145 x145 xm145 1.51094605540703e-12
Vx145 xm145 0 0
Gx145_2 x145 0 u2 0 -0.0541338253751461
Rx146 x146 0 1
Fxc146_145 x146 0 Vx145 -1.32367213232931
Cx146 x146 xm146 1.51094605540703e-12
Vx146 xm146 0 0
Gx146_2 x146 0 u2 0 0.071655436065462
Rx147 x147 0 1
Fxc147_148 x147 0 Vx148 26.4827669935933
Cx147 x147 xm147 1.70972884859627e-12
Vx147 xm147 0 0
Gx147_2 x147 0 u2 0 -0.0157240174750674
Rx148 x148 0 1
Fxc148_147 x148 0 Vx147 -3.41762555710375
Cx148 x148 xm148 1.70972884859627e-12
Vx148 xm148 0 0
Gx148_2 x148 0 u2 0 0.0537388039831365
Rx149 x149 0 1
Fxc149_150 x149 0 Vx150 4.90806690144271
Cx149 x149 xm149 1.61515298397391e-12
Vx149 xm149 0 0
Gx149_2 x149 0 u2 0 -0.0053071238425388
Rx150 x150 0 1
Fxc150_149 x150 0 Vx149 -31.8385219732171
Cx150 x150 xm150 1.61515298397391e-12
Vx150 xm150 0 0
Gx150_2 x150 0 u2 0 0.168970979075256
Rx151 x151 0 1
Fxc151_152 x151 0 Vx152 3.33564145012427
Cx151 x151 xm151 3.3832600882424e-12
Vx151 xm151 0 0
Gx151_2 x151 0 u2 0 -0.107401191029852
Rx152 x152 0 1
Fxc152_151 x152 0 Vx151 -10.4705516268112
Cx152 x152 xm152 3.3832600882424e-12
Vx152 xm152 0 0
Gx152_2 x152 0 u2 0 1.12454971545908
Rx153 x153 0 1
Fxc153_154 x153 0 Vx154 4.59607910724032
Cx153 x153 xm153 6.36249392361281e-12
Vx153 xm153 0 0
Gx153_2 x153 0 u2 0 -0.219549995998787
Rx154 x154 0 1
Fxc154_153 x154 0 Vx153 -3.70326767108602
Cx154 x154 xm154 6.36249392361281e-12
Vx154 xm154 0 0
Gx154_2 x154 0 u2 0 0.813052402369373
Rx155 x155 0 1
Fxc155_156 x155 0 Vx156 31.1087663218418
Cx155 x155 xm155 4.08890323417608e-12
Vx155 xm155 0 0
Gx155_2 x155 0 u2 0 -0.00446614223321578
Rx156 x156 0 1
Fxc156_155 x156 0 Vx155 -1.71066564091351
Cx156 x156 xm156 4.08890323417608e-12
Vx156 xm156 0 0
Gx156_2 x156 0 u2 0 0.00764007606579495
Rx157 x157 0 1
Fxc157_158 x157 0 Vx158 5.71439220701276
Cx157 x157 xm157 1.41898003518717e-11
Vx157 xm157 0 0
Gx157_2 x157 0 u2 0 -0.560700405408673
Rx158 x158 0 1
Fxc158_157 x158 0 Vx157 -1.16884670902194
Cx158 x158 xm158 1.41898003518717e-11
Vx158 xm158 0 0
Gx158_2 x158 0 u2 0 0.655372823609195
Rx159 x159 0 1
Fxc159_160 x159 0 Vx160 1.72311443495368
Cx159 x159 xm159 3.02223658791127e-11
Vx159 xm159 0 0
Gx159_2 x159 0 u2 0 -0.628812427346403
Rx160 x160 0 1
Fxc160_159 x160 0 Vx159 -1.42723657161402
Cx160 x160 xm160 3.02223658791127e-11
Vx160 xm160 0 0
Gx160_2 x160 0 u2 0 0.897464092994171
Rx161 x161 0 1
Fxc161_162 x161 0 Vx162 3.90044888591569
Cx161 x161 xm161 1.30273315544064e-11
Vx161 xm161 0 0
Gx161_2 x161 0 u2 0 -0.00042427500476389
Rx162 x162 0 1
Fxc162_161 x162 0 Vx161 -7.64492386011162
Cx162 x162 xm162 1.30273315544064e-11
Vx162 xm162 0 0
Gx162_2 x162 0 u2 0 0.00324355010716844
Rx163 x163 0 1
Fxc163_164 x163 0 Vx164 14.6886133860057
Cx163 x163 xm163 4.87133831260231e-12
Vx163 xm163 0 0
Gx163_2 x163 0 u2 0 -2.337291065694e-05
Rx164 x164 0 1
Fxc164_163 x164 0 Vx163 -18.5859597307902
Cx164 x164 xm164 4.87133831260231e-12
Vx164 xm164 0 0
Gx164_2 x164 0 u2 0 0.000434407976261244
Rx165 x165 0 1
Fxc165_166 x165 0 Vx166 0.883423787931558
Cx165 x165 xm165 7.06557064659634e-11
Vx165 xm165 0 0
Gx165_2 x165 0 u2 0 -0.153494392321192
Rx166 x166 0 1
Fxc166_165 x166 0 Vx165 -1.70926725354214
Cx166 x166 xm166 7.06557064659634e-11
Vx166 xm166 0 0
Gx166_2 x166 0 u2 0 0.262362938396962
Rx167 x167 0 1
Fxc167_168 x167 0 Vx168 124.098488416375
Cx167 x167 xm167 9.00586691578378e-12
Vx167 xm167 0 0
Gx167_2 x167 0 u2 0 -1.47921737094881e-05
Rx168 x168 0 1
Fxc168_167 x168 0 Vx167 -2.75761814643032
Cx168 x168 xm168 9.00586691578378e-12
Vx168 xm168 0 0
Gx168_2 x168 0 u2 0 4.0791166646434e-05
Rx169 x169 0 1
Fxc169_170 x169 0 Vx170 163.851006608003
Cx169 x169 xm169 6.72924348226814e-13
Vx169 xm169 0 0
Gx169_2 x169 0 u2 0 -1.57729814895469e-08
Rx170 x170 0 1
Fxc170_169 x170 0 Vx169 -387.360098261158
Cx170 x170 xm170 6.72924348226814e-13
Vx170 xm170 0 0
Gx170_2 x170 0 u2 0 6.10982365966232e-06
Rx171 x171 0 1
Fxc171_172 x171 0 Vx172 306.207387820098
Cx171 x171 xm171 7.40586010206479e-13
Vx171 xm171 0 0
Gx171_2 x171 0 u2 0 -2.41648663461334e-08
Rx172 x172 0 1
Fxc172_171 x172 0 Vx171 -194.551709607962
Cx172 x172 xm172 7.40586010206479e-13
Vx172 xm172 0 0
Gx172_2 x172 0 u2 0 4.70131606008815e-06
Rx173 x173 0 1
Fxc173_174 x173 0 Vx174 0.0160355726388108
Cx173 x173 xm173 2.7189670410967e-10
Vx173 xm173 0 0
Gx173_2 x173 0 u2 0 -0.252181174893651
Rx174 x174 0 1
Fxc174_173 x174 0 Vx173 -0.385129907307044
Cx174 x174 xm174 2.7189670410967e-10
Vx174 xm174 0 0
Gx174_2 x174 0 u2 0 0.0971225125113733
Rx175 x175 0 1
Fxc175_176 x175 0 Vx176 3883.8368971596
Cx175 x175 xm175 3.4033679671408e-13
Vx175 xm175 0 0
Gx175_2 x175 0 u2 0 -6.43742142732494e-09
Rx176 x176 0 1
Fxc176_175 x176 0 Vx175 -83.2679881232261
Cx176 x176 xm176 3.40336796714079e-13
Vx176 xm176 0 0
Gx176_2 x176 0 u2 0 5.36031130954695e-07
Rx177 x177 0 1
Fxc177_178 x177 0 Vx178 5.0724427210576
Cx177 x177 xm177 1.77838009044698e-11
Vx177 xm177 0 0
Gx177_2 x177 0 u2 0 -6.61619443070564e-05
Rx178 x178 0 1
Fxc178_177 x178 0 Vx177 -25.0008412330546
Cx178 x178 xm178 1.77838009044698e-11
Vx178 xm178 0 0
Gx178_2 x178 0 u2 0 0.00165410426529092
Rx179 x179 0 1
Fxc179_180 x179 0 Vx180 13845.9175377635
Cx179 x179 xm179 6.45459166206642e-14
Vx179 xm179 0 0
Gx179_2 x179 0 u2 0 -1.69814103132952e-09
Rx180 x180 0 1
Fxc180_179 x180 0 Vx179 -725.195731764376
Cx180 x180 xm180 6.45459166206643e-14
Vx180 xm180 0 0
Gx180_2 x180 0 u2 0 1.23148462785412e-06
Rx181 x181 0 1
Fxc181_182 x181 0 Vx182 39.6679773982074
Cx181 x181 xm181 3.60587813907164e-12
Vx181 xm181 0 0
Gx181_2 x181 0 u2 0 -7.30635638620476e-07
Rx182 x182 0 1
Fxc182_181 x182 0 Vx181 -85.5570048481699
Cx182 x182 xm182 3.60587813907164e-12
Vx182 xm182 0 0
Gx182_2 x182 0 u2 0 6.25109968756977e-05
Rx183 x183 0 1
Fxc183_184 x183 0 Vx184 17.5544024554666
Cx183 x183 xm183 1.33799391561211e-11
Vx183 xm183 0 0
Gx183_2 x183 0 u2 0 -6.30271842872257e-05
Rx184 x184 0 1
Fxc184_183 x184 0 Vx183 -16.22048460148
Cx184 x184 xm184 1.33799391561211e-11
Vx184 xm184 0 0
Gx184_2 x184 0 u2 0 0.00102233147220559
Rx185 x185 0 1
Fxc185_186 x185 0 Vx186 6.47967426392752
Cx185 x185 xm185 2.86431819527606e-12
Vx185 xm185 0 0
Gx185_2 x185 0 u2 0 -5.60577663614379e-08
Rx186 x186 0 1
Fxc186_185 x186 0 Vx185 -892.679963091082
Cx186 x186 xm186 2.86431819527606e-12
Vx186 xm186 0 0
Gx186_2 x186 0 u2 0 5.00416448064969e-05
Rx187 x187 0 1
Fxc187_188 x187 0 Vx188 16.3853652031555
Cx187 x187 xm187 7.0808537117008e-12
Vx187 xm187 0 0
Gx187_2 x187 0 u2 0 -4.08177704341213e-06
Rx188 x188 0 1
Fxc188_187 x188 0 Vx187 -65.7192053528268
Cx188 x188 xm188 7.0808537117008e-12
Vx188 xm188 0 0
Gx188_2 x188 0 u2 0 0.000268251143720456
Rx189 x189 0 1
Fxc189_190 x189 0 Vx190 191.492139995185
Cx189 x189 xm189 8.39484573603046e-12
Vx189 xm189 0 0
Gx189_2 x189 0 u2 0 -6.84059839155567e-06
Rx190 x190 0 1
Fxc190_189 x190 0 Vx189 -4.51660616312773
Cx190 x190 xm190 8.39484573603046e-12
Vx190 xm190 0 0
Gx190_2 x190 0 u2 0 3.0896288854782e-05
Rx191 x191 0 1
Fxc191_192 x191 0 Vx192 1656.04860406475
Cx191 x191 xm191 2.83045279415423e-13
Vx191 xm191 0 0
Gx191_2 x191 0 u2 0 -5.52656520350403e-09
Rx192 x192 0 1
Fxc192_191 x192 0 Vx191 -483.660340290366
Cx192 x192 xm192 2.83045279415423e-13
Vx192 xm192 0 0
Gx192_2 x192 0 u2 0 2.67298040696365e-06
Rx193 x193 0 1
Fxc193_194 x193 0 Vx194 28.4254838316825
Cx193 x193 xm193 5.19274272676225e-12
Vx193 xm193 0 0
Gx193_2 x193 0 u2 0 -4.9669277694326e-07
Rx194 x194 0 1
Fxc194_193 x194 0 Vx193 -94.7959216516197
Cx194 x194 xm194 5.19274272676225e-12
Vx194 xm194 0 0
Gx194_2 x194 0 u2 0 4.70844495680387e-05
Rx195 x195 0 1
Fxc195_196 x195 0 Vx196 1486.56318758971
Cx195 x195 xm195 6.76962091359381e-13
Vx195 xm195 0 0
Gx195_2 x195 0 u2 0 -3.76801335160697e-09
Rx196 x196 0 1
Fxc196_195 x196 0 Vx195 -115.571696649177
Cx196 x196 xm196 6.76962091359381e-13
Vx196 xm196 0 0
Gx196_2 x196 0 u2 0 4.3547569604197e-07
Rx197 x197 0 1
Fxc197_198 x197 0 Vx198 8.04710451777268
Cx197 x197 xm197 1.60390660485385e-11
Vx197 xm197 0 0
Gx197_2 x197 0 u2 0 -1.32944560028944e-05
Rx198 x198 0 1
Fxc198_197 x198 0 Vx197 -39.1667918819358
Cx198 x198 xm198 1.60390660485385e-11
Vx198 xm198 0 0
Gx198_2 x198 0 u2 0 0.000520701191448915
Rx199 x199 0 1
Fxc199_200 x199 0 Vx200 12.5358545634304
Cx199 x199 xm199 3.65373015413682e-11
Vx199 xm199 0 0
Gx199_2 x199 0 u2 0 -0.0001364299139217
Rx200 x200 0 1
Fxc200_199 x200 0 Vx199 -5.52335113139414
Cx200 x200 xm200 3.65373015413682e-11
Vx200 xm200 0 0
Gx200_2 x200 0 u2 0 0.000753550319415429
Rx201 x201 0 1
Fxc201_202 x201 0 Vx202 182.671903429941
Cx201 x201 xm201 4.9605444448296e-12
Vx201 xm201 0 0
Gx201_2 x201 0 u2 0 -4.08322597091157e-07
Rx202 x202 0 1
Fxc202_201 x202 0 Vx201 -25.1794023490687
Cx202 x202 xm202 4.9605444448296e-12
Vx202 xm202 0 0
Gx202_2 x202 0 u2 0 1.02813189603749e-05
Rx203 x203 0 1
Fxc203_204 x203 0 Vx204 2319.34205346775
Cx203 x203 xm203 1.85213203877505e-12
Vx203 xm203 0 0
Gx203_2 x203 0 u2 0 -7.69925061565872e-08
Rx204 x204 0 1
Fxc204_203 x204 0 Vx203 -15.8696730598753
Cx204 x204 xm204 1.85213203877505e-12
Vx204 xm204 0 0
Gx204_2 x204 0 u2 0 1.22184590076548e-06
Rx205 x205 0 1
Fxc205_206 x205 0 Vx206 19.3941995504026
Cx205 x205 xm205 6.12244434678794e-12
Vx205 xm205 0 0
Gx205_2 x205 0 u2 0 -1.24322943943029e-07
Rx206 x206 0 1
Fxc206_205 x206 0 Vx205 -203.052911765391
Cx206 x206 xm206 6.12244434678794e-12
Vx206 xm206 0 0
Gx206_2 x206 0 u2 0 2.52441357668775e-05
Rx207 x207 0 1
Fxc207_208 x207 0 Vx208 279.030231190825
Cx207 x207 xm207 1.14029529690273e-12
Vx207 xm207 0 0
Gx207_2 x207 0 u2 0 -1.48115637776197e-08
Rx208 x208 0 1
Fxc208_207 x208 0 Vx207 -469.564820772117
Cx208 x208 xm208 1.14029529690273e-12
Vx208 xm208 0 0
Gx208_2 x208 0 u2 0 6.95498929059279e-06
Rx209 x209 0 1
Fxc209_210 x209 0 Vx210 18.7137522961697
Cx209 x209 xm209 9.47069571391727e-12
Vx209 xm209 0 0
Gx209_2 x209 0 u2 0 -3.46891155417485e-07
Rx210 x210 0 1
Fxc210_209 x210 0 Vx209 -113.001417510361
Cx210 x210 xm210 9.47069571391727e-12
Vx210 xm210 0 0
Gx210_2 x210 0 u2 0 3.91991922839827e-05
Rx211 x211 0 1
Fxc211_212 x211 0 Vx212 479.227528848619
Cx211 x211 xm211 1.41828331495617e-12
Vx211 xm211 0 0
Gx211_2 x211 0 u2 0 -3.08696535426107e-08
Rx212 x212 0 1
Fxc212_211 x212 0 Vx211 -211.377370000322
Cx212 x212 xm212 1.41828331495617e-12
Vx212 xm212 0 0
Gx212_2 x212 0 u2 0 6.52514617865817e-06
Rx213 x213 0 1
Fxc213_214 x213 0 Vx214 78.1405959847492
Cx213 x213 xm213 5.0878616870562e-12
Vx213 xm213 0 0
Gx213_2 x213 0 u2 0 -6.25008907744157e-08
Rx214 x214 0 1
Fxc214_213 x214 0 Vx213 -121.608587323861
Cx214 x214 xm214 5.0878616870562e-12
Vx214 xm214 0 0
Gx214_2 x214 0 u2 0 7.60064503355961e-06
Rx215 x215 0 1
Fxc215_216 x215 0 Vx216 14.4409176695634
Cx215 x215 xm215 4.66368852903178e-11
Vx215 xm215 0 0
Gx215_2 x215 0 u2 0 -1.63588376035471e-05
Rx216 x216 0 1
Fxc216_215 x216 0 Vx215 -10.1072334903951
Cx216 x216 xm216 4.66368852903178e-11
Vx216 xm216 0 0
Gx216_2 x216 0 u2 0 0.000165342591290507
Rx217 x217 0 1
Fxc217_218 x217 0 Vx218 24.9417241299353
Cx217 x217 xm217 5.38073810888037e-12
Vx217 xm217 0 0
Gx217_2 x217 0 u2 0 -4.0176242497223e-08
Rx218 x218 0 1
Fxc218_217 x218 0 Vx217 -391.968506784494
Cx218 x218 xm218 5.38073810888037e-12
Vx218 xm218 0 0
Gx218_2 x218 0 u2 0 1.57478217798482e-05
Rx219 x219 0 1
Fxc219_220 x219 0 Vx220 32.3912574676233
Cx219 x219 xm219 9.45572193374133e-12
Vx219 xm219 0 0
Gx219_2 x219 0 u2 0 -3.2730727813511e-07
Rx220 x220 0 1
Fxc220_219 x220 0 Vx219 -123.785718346195
Cx220 x220 xm220 9.45572193374133e-12
Vx220 xm220 0 0
Gx220_2 x220 0 u2 0 4.05159665438925e-05
Rx221 x221 0 1
Fxc221_222 x221 0 Vx222 121.441340165187
Cx221 x221 xm221 1.20602139754355e-11
Vx221 xm221 0 0
Gx221_2 x221 0 u2 0 -2.80614515104026e-07
Rx222 x222 0 1
Fxc222_221 x222 0 Vx221 -24.3479652283957
Cx222 x222 xm222 1.20602139754355e-11
Vx222 xm222 0 0
Gx222_2 x222 0 u2 0 6.83239245633593e-06
Rx223 x223 0 1
Fxc223_224 x223 0 Vx224 49.6168852878725
Cx223 x223 xm223 1.25498339510922e-11
Vx223 xm223 0 0
Gx223_2 x223 0 u2 0 -1.95746963053652e-07
Rx224 x224 0 1
Fxc224_223 x224 0 Vx223 -75.9764171568511
Cx224 x224 xm224 1.25498339510922e-11
Vx224 xm224 0 0
Gx224_2 x224 0 u2 0 1.4872152922151e-05
Rx225 x225 0 1
Fxc225_226 x225 0 Vx226 63.8706653122786
Cx225 x225 xm225 3.32631261202093e-11
Vx225 xm225 0 0
Gx225_2 x225 0 u2 0 -1.49792822621642e-06
Rx226 x226 0 1
Fxc226_225 x226 0 Vx225 -14.84313463802
Cx226 x226 xm226 3.32631261202093e-11
Vx226 xm226 0 0
Gx226_2 x226 0 u2 0 2.22339503398209e-05
Rx227 x227 0 1
Fxc227_228 x227 0 Vx228 12.031017822058
Cx227 x227 xm227 1.45379770932265e-10
Vx227 xm227 0 0
Gx227_2 x227 0 u2 0 -4.96721675520996e-05
Rx228 x228 0 1
Fxc228_227 x228 0 Vx227 -5.44480279773338
Cx228 x228 xm228 1.45379770932265e-10
Vx228 xm228 0 0
Gx228_2 x228 0 u2 0 0.000270455156857153
Rx229 x229 0 1
Fxc229_230 x229 0 Vx230 2.9714146688483
Cx229 x229 xm229 4.64722716786655e-11
Vx229 xm229 0 0
Gx229_2 x229 0 u2 0 -3.08955271269557e-07
Rx230 x230 0 1
Fxc230_229 x230 0 Vx229 -1104.36334765002
Cx230 x230 xm230 4.64722716786655e-11
Vx230 xm230 0 0
Gx230_2 x230 0 u2 0 0.000341198877653368
Rx231 x231 0 1
Fxc231_232 x231 0 Vx232 5.20140854675853
Cx231 x231 xm231 2.59641851055736e-10
Vx231 xm231 0 0
Gx231_2 x231 0 u2 0 -8.29583888406763e-06
Rx232 x232 0 1
Fxc232_231 x232 0 Vx231 -91.2119786642537
Cx232 x232 xm232 2.59641851055736e-10
Vx232 xm232 0 0
Gx232_2 x232 0 u2 0 0.000756679879295663
Rx233 x233 0 1
Fxc233_234 x233 0 Vx234 0.062263861302183
Cx233 x233 xm233 6.69011915274045e-09
Vx233 xm233 0 0
Gx233_2 x233 0 u2 0 -0.00132873780325519
Rx234 x234 0 1
Fxc234_233 x234 0 Vx233 -80.1316415743038
Cx234 x234 xm234 6.69011915274045e-09
Vx234 xm234 0 0
Gx234_2 x234 0 u2 0 0.106473941396673
Rx235 x235 0 1
Fxc235_236 x235 0 Vx236 0.548055024070288
Cx235 x235 xm235 1.52744488718003e-09
Vx235 xm235 0 0
Gx235_2 x235 0 u2 0 -7.37971537747601e-05
Rx236 x236 0 1
Fxc236_235 x236 0 Vx235 -53.639435375902
Cx236 x236 xm236 1.52744488718003e-09
Vx236 xm236 0 0
Gx236_2 x236 0 u2 0 0.00395843766082675
Rx237 x237 0 1
Fxc237_238 x237 0 Vx238 340.632664606375
Cx237 x237 xm237 1.70618985523348e-11
Vx237 xm237 0 0
Gx237_2 x237 0 u2 0 -1.21812298740389e-06
Rx238 x238 0 1
Fxc238_237 x238 0 Vx237 -102.367409115388
Cx238 x238 xm238 1.70618985523348e-11
Vx238 xm238 0 0
Gx238_2 x238 0 u2 0 0.000124696094204433
Rx239 x239 0 1
Cx239 x239 0 1.12913277439532e-08
Gx239_2 x239 0 u2 0 -0.962863269901288
Rx240 x240 0 1
Cx240 x240 0 2.13606987450335e-08
Gx240_2 x240 0 u2 0 -1.07499798049592
Gyc1_1 y1 0 x1 0 0.476755492360765
Gyc1_2 y1 0 x2 0 1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 0.743068576843484
Gyc1_5 y1 0 x5 0 1
Gyc1_6 y1 0 x6 0 -0.041213958771277
Gyc1_7 y1 0 x7 0 1
Gyc1_8 y1 0 x8 0 -1
Gyc1_9 y1 0 x9 0 0.833953803673922
Gyc1_10 y1 0 x10 0 -0.0920525661127817
Gyc1_11 y1 0 x11 0 0.341495855032085
Gyc1_12 y1 0 x12 0 -0.347439715194234
Gyc1_13 y1 0 x13 0 -0.19329456952945
Gyc1_14 y1 0 x14 0 1
Gyc1_15 y1 0 x15 0 -1
Gyc1_16 y1 0 x16 0 -1
Gyc1_17 y1 0 x17 0 0.189970478779657
Gyc1_18 y1 0 x18 0 -1
Gyc1_19 y1 0 x19 0 1
Gyc1_20 y1 0 x20 0 -0.172229036544693
Gyc1_21 y1 0 x21 0 -0.0111836591709204
Gyc1_22 y1 0 x22 0 -0.868471803499502
Gyc1_23 y1 0 x23 0 0.0384169549193403
Gyc1_24 y1 0 x24 0 -1
Gyc1_25 y1 0 x25 0 -1
Gyc1_26 y1 0 x26 0 -1
Gyc1_27 y1 0 x27 0 1
Gyc1_28 y1 0 x28 0 -1
Gyc1_29 y1 0 x29 0 -0.883701549728683
Gyc1_30 y1 0 x30 0 0.606126734097666
Gyc1_31 y1 0 x31 0 -0.684282210886985
Gyc1_32 y1 0 x32 0 -1
Gyc1_33 y1 0 x33 0 -0.847792853556691
Gyc1_34 y1 0 x34 0 0.336463903482262
Gyc1_35 y1 0 x35 0 0.0693513462455304
Gyc1_36 y1 0 x36 0 0.0769430454579666
Gyc1_37 y1 0 x37 0 0.96668125244406
Gyc1_38 y1 0 x38 0 0.279440230917415
Gyc1_39 y1 0 x39 0 -0.991068612783289
Gyc1_40 y1 0 x40 0 -1
Gyc1_41 y1 0 x41 0 -0.422500097856906
Gyc1_42 y1 0 x42 0 0.535554728817061
Gyc1_43 y1 0 x43 0 0.27669789824258
Gyc1_44 y1 0 x44 0 0.342654436373517
Gyc1_45 y1 0 x45 0 -0.00589668033550414
Gyc1_46 y1 0 x46 0 -0.592821144154977
Gyc1_47 y1 0 x47 0 0.14964604391448
Gyc1_48 y1 0 x48 0 -0.0858723840751985
Gyc1_49 y1 0 x49 0 -0.0823703862530285
Gyc1_50 y1 0 x50 0 0.0593893489872369
Gyc1_51 y1 0 x51 0 1
Gyc1_52 y1 0 x52 0 -0.0656042776603331
Gyc1_53 y1 0 x53 0 -0.056529171908485
Gyc1_54 y1 0 x54 0 0.0939675143721512
Gyc1_55 y1 0 x55 0 -0.131192317209834
Gyc1_56 y1 0 x56 0 0.0290052661857464
Gyc1_57 y1 0 x57 0 -0.058876875355895
Gyc1_58 y1 0 x58 0 -0.0575405943986204
Gyc1_59 y1 0 x59 0 0.172724898134539
Gyc1_60 y1 0 x60 0 -0.0207300139029315
Gyc1_61 y1 0 x61 0 0.0835482483816108
Gyc1_62 y1 0 x62 0 -0.0414053830932768
Gyc1_63 y1 0 x63 0 0.363923183598804
Gyc1_64 y1 0 x64 0 -0.0435734133268087
Gyc1_65 y1 0 x65 0 0.0674474538144532
Gyc1_66 y1 0 x66 0 0.0103492442132175
Gyc1_67 y1 0 x67 0 -0.0416532742332278
Gyc1_68 y1 0 x68 0 -0.0109825064449007
Gyc1_69 y1 0 x69 0 -0.0156125127162462
Gyc1_70 y1 0 x70 0 -0.0554656434441262
Gyc1_71 y1 0 x71 0 0.0472612189646481
Gyc1_72 y1 0 x72 0 -0.0882719285640275
Gyc1_73 y1 0 x73 0 0.0108200873040445
Gyc1_74 y1 0 x74 0 0.0797566489755668
Gyc1_75 y1 0 x75 0 0.125380852357917
Gyc1_76 y1 0 x76 0 0.0409941195742907
Gyc1_77 y1 0 x77 0 -0.0106304845527899
Gyc1_78 y1 0 x78 0 0.232643223743051
Gyc1_79 y1 0 x79 0 0.65284506613295
Gyc1_80 y1 0 x80 0 -0.0255628708183149
Gyc1_81 y1 0 x81 0 0.0556254105132815
Gyc1_82 y1 0 x82 0 -0.115918325897544
Gyc1_83 y1 0 x83 0 0.467424356798958
Gyc1_84 y1 0 x84 0 -0.0745346105151354
Gyc1_85 y1 0 x85 0 0.040364583950051
Gyc1_86 y1 0 x86 0 -0.0316955648736634
Gyc1_87 y1 0 x87 0 -0.0948599338059692
Gyc1_88 y1 0 x88 0 0.239142197714386
Gyc1_89 y1 0 x89 0 0.007641802372743
Gyc1_90 y1 0 x90 0 0.477329488314415
Gyc1_91 y1 0 x91 0 0.056948119702977
Gyc1_92 y1 0 x92 0 0.000869017318908231
Gyc1_93 y1 0 x93 0 -0.0271763116165014
Gyc1_94 y1 0 x94 0 0.00666888461765092
Gyc1_95 y1 0 x95 0 -0.0224373052838726
Gyc1_96 y1 0 x96 0 0.00255237868733906
Gyc1_97 y1 0 x97 0 -0.0431001185910109
Gyc1_98 y1 0 x98 0 -0.0273575251072095
Gyc1_99 y1 0 x99 0 0.00517649547116734
Gyc1_100 y1 0 x100 0 0.00352539508714368
Gyc1_101 y1 0 x101 0 -0.010719137178815
Gyc1_102 y1 0 x102 0 -0.0164402423140159
Gyc1_103 y1 0 x103 0 0.00702114408848533
Gyc1_104 y1 0 x104 0 -0.0306766597498111
Gyc1_105 y1 0 x105 0 0.0253102031282351
Gyc1_106 y1 0 x106 0 0.0713232186971717
Gyc1_107 y1 0 x107 0 0.0261962924935928
Gyc1_108 y1 0 x108 0 -0.0463478036819396
Gyc1_109 y1 0 x109 0 0.0457264458408878
Gyc1_110 y1 0 x110 0 0.243395047311055
Gyc1_111 y1 0 x111 0 -0.0187979939078364
Gyc1_112 y1 0 x112 0 -0.0378046409991195
Gyc1_113 y1 0 x113 0 0.00331396542485066
Gyc1_114 y1 0 x114 0 -0.00401043740348861
Gyc1_115 y1 0 x115 0 -0.0861893125965617
Gyc1_116 y1 0 x116 0 -0.00213149387720721
Gyc1_117 y1 0 x117 0 -0.0635537292098876
Gyc1_118 y1 0 x118 0 -0.12729274009847
Gyc1_119 y1 0 x119 0 -0.935341016212936
Gyc1_120 y1 0 x120 0 0.0077718245969283
Gyc1_121 y1 0 x121 0 0.170570259702434
Gyc1_122 y1 0 x122 0 -0.322402002415916
Gyc1_123 y1 0 x123 0 -0.362381754874188
Gyc1_124 y1 0 x124 0 0.0260863247614053
Gyc1_125 y1 0 x125 0 -0.16528432280057
Gyc1_126 y1 0 x126 0 0.757468656084447
Gyc1_127 y1 0 x127 0 -0.809850468895608
Gyc1_128 y1 0 x128 0 -0.0498644578897116
Gyc1_129 y1 0 x129 0 0.220683291074479
Gyc1_130 y1 0 x130 0 -0.296072896536621
Gyc1_131 y1 0 x131 0 -0.359250994759376
Gyc1_132 y1 0 x132 0 -0.257175169091255
Gyc1_133 y1 0 x133 0 -1
Gyc1_134 y1 0 x134 0 -0.0841563217810921
Gyc1_135 y1 0 x135 0 -0.590216795928101
Gyc1_136 y1 0 x136 0 0.394429943095389
Gyc1_137 y1 0 x137 0 0.47494755111382
Gyc1_138 y1 0 x138 0 0.879382258459141
Gyc1_139 y1 0 x139 0 0.202339479098439
Gyc1_140 y1 0 x140 0 0.669704528793534
Gyc1_141 y1 0 x141 0 -0.266127141981907
Gyc1_142 y1 0 x142 0 -0.0535307167887532
Gyc1_143 y1 0 x143 0 0.625327720773989
Gyc1_144 y1 0 x144 0 -0.12938804235411
Gyc1_145 y1 0 x145 0 -0.28429544191859
Gyc1_146 y1 0 x146 0 0.00900995582973229
Gyc1_147 y1 0 x147 0 -0.468867765984496
Gyc1_148 y1 0 x148 0 0.145444736955072
Gyc1_149 y1 0 x149 0 -0.53147171173106
Gyc1_150 y1 0 x150 0 -0.144073229610815
Gyc1_151 y1 0 x151 0 0.220707090235644
Gyc1_152 y1 0 x152 0 0.309471466626329
Gyc1_153 y1 0 x153 0 0.360727833674599
Gyc1_154 y1 0 x154 0 -0.267122271181811
Gyc1_155 y1 0 x155 0 0.108662479376099
Gyc1_156 y1 0 x156 0 -0.987053463594075
Gyc1_157 y1 0 x157 0 -0.230456416951238
Gyc1_158 y1 0 x158 0 -0.150920137989355
Gyc1_159 y1 0 x159 0 0.242101615189885
Gyc1_160 y1 0 x160 0 0.0931044340476121
Gyc1_161 y1 0 x161 0 -0.462212611330448
Gyc1_162 y1 0 x162 0 0.145930727549391
Gyc1_163 y1 0 x163 0 0.117162057880996
Gyc1_164 y1 0 x164 0 0.1573883553426
Gyc1_165 y1 0 x165 0 -0.239948038884739
Gyc1_166 y1 0 x166 0 -0.0346387253870144
Gyc1_167 y1 0 x167 0 -0.2858653331517
Gyc1_168 y1 0 x168 0 -0.303652395482837
Gyc1_169 y1 0 x169 0 0.290909940553729
Gyc1_170 y1 0 x170 0 0.272075308264826
Gyc1_171 y1 0 x171 0 -0.300022994813327
Gyc1_172 y1 0 x172 0 -0.17117234642604
Gyc1_173 y1 0 x173 0 -0.152518541644732
Gyc1_174 y1 0 x174 0 -0.151900884747415
Gyc1_175 y1 0 x175 0 0.257781194959736
Gyc1_176 y1 0 x176 0 0.246242315105429
Gyc1_177 y1 0 x177 0 -0.0653598301113363
Gyc1_178 y1 0 x178 0 -0.234355951088827
Gyc1_179 y1 0 x179 0 -0.00298398632806263
Gyc1_180 y1 0 x180 0 -0.137509383320347
Gyc1_181 y1 0 x181 0 -0.358540704732373
Gyc1_182 y1 0 x182 0 -0.236409859087956
Gyc1_183 y1 0 x183 0 -0.36128830453544
Gyc1_184 y1 0 x184 0 -0.192500403801402
Gyc1_185 y1 0 x185 0 -0.472215514040229
Gyc1_186 y1 0 x186 0 -0.290254313003358
Gyc1_187 y1 0 x187 0 -0.106905403055082
Gyc1_188 y1 0 x188 0 0.332477314335591
Gyc1_189 y1 0 x189 0 -0.283517162262608
Gyc1_190 y1 0 x190 0 0.874040828075563
Gyc1_191 y1 0 x191 0 0.0236440810725644
Gyc1_192 y1 0 x192 0 0.212037147520515
Gyc1_193 y1 0 x193 0 0.0260055879151504
Gyc1_194 y1 0 x194 0 -0.401729221411483
Gyc1_195 y1 0 x195 0 1
Gyc1_196 y1 0 x196 0 -0.434946355661435
Gyc1_197 y1 0 x197 0 -0.167004509391515
Gyc1_198 y1 0 x198 0 -0.307010291386517
Gyc1_199 y1 0 x199 0 -0.407577870763658
Gyc1_200 y1 0 x200 0 -0.0613548038805823
Gyc1_201 y1 0 x201 0 -0.167753015862616
Gyc1_202 y1 0 x202 0 0.666328117718069
Gyc1_203 y1 0 x203 0 -0.168362745210874
Gyc1_204 y1 0 x204 0 1
Gyc1_205 y1 0 x205 0 -0.754797227992288
Gyc1_206 y1 0 x206 0 -0.191960779011339
Gyc1_207 y1 0 x207 0 0.00771586718421072
Gyc1_208 y1 0 x208 0 -0.138822252704161
Gyc1_209 y1 0 x209 0 0.26534263116608
Gyc1_210 y1 0 x210 0 -0.288937935797905
Gyc1_211 y1 0 x211 0 -0.0134864164905471
Gyc1_212 y1 0 x212 0 -0.290630899856317
Gyc1_213 y1 0 x213 0 0.69971041223303
Gyc1_214 y1 0 x214 0 0.0287794389404482
Gyc1_215 y1 0 x215 0 0.45701767435967
Gyc1_216 y1 0 x216 0 -0.144003983164729
Gyc1_217 y1 0 x217 0 0.49021210906903
Gyc1_218 y1 0 x218 0 0.211412346826374
Gyc1_219 y1 0 x219 0 -0.141887832821391
Gyc1_220 y1 0 x220 0 -0.218588424785986
Gyc1_221 y1 0 x221 0 0.304321033209898
Gyc1_222 y1 0 x222 0 -1
Gyc1_223 y1 0 x223 0 0.513684100825841
Gyc1_224 y1 0 x224 0 0.0499001028095081
Gyc1_225 y1 0 x225 0 -0.17014920064632
Gyc1_226 y1 0 x226 0 0.564058475348216
Gyc1_227 y1 0 x227 0 0.0557675892264094
Gyc1_228 y1 0 x228 0 0.334452732436301
Gyc1_229 y1 0 x229 0 -0.527778555517625
Gyc1_230 y1 0 x230 0 0.047554287508261
Gyc1_231 y1 0 x231 0 0.0868227501259418
Gyc1_232 y1 0 x232 0 0.00759524125061287
Gyc1_233 y1 0 x233 0 0.549227837438885
Gyc1_234 y1 0 x234 0 -0.0162927261691346
Gyc1_235 y1 0 x235 0 0.104673391300026
Gyc1_236 y1 0 x236 0 -0.032323803006195
Gyc1_237 y1 0 x237 0 -0.0527646552617197
Gyc1_238 y1 0 x238 0 -0.0131194778952336
Gyc1_239 y1 0 x239 0 0.0683838858236863
Gyc1_240 y1 0 x240 0 -0.02924420805896
Gyc2_1 y2 0 x1 0 1
Gyc2_2 y2 0 x2 0 0.16762580141293
Gyc2_3 y2 0 x3 0 -0.361758137944807
Gyc2_4 y2 0 x4 0 1
Gyc2_5 y2 0 x5 0 -0.380163459903739
Gyc2_6 y2 0 x6 0 1
Gyc2_7 y2 0 x7 0 0.201798184789728
Gyc2_8 y2 0 x8 0 0.257867242752703
Gyc2_9 y2 0 x9 0 1
Gyc2_10 y2 0 x10 0 1
Gyc2_11 y2 0 x11 0 1
Gyc2_12 y2 0 x12 0 -1
Gyc2_13 y2 0 x13 0 1
Gyc2_14 y2 0 x14 0 -0.632080101007903
Gyc2_15 y2 0 x15 0 0.290486823149051
Gyc2_16 y2 0 x16 0 0.0697994475542055
Gyc2_17 y2 0 x17 0 1
Gyc2_18 y2 0 x18 0 0.0210736921059279
Gyc2_19 y2 0 x19 0 0.903615554375801
Gyc2_20 y2 0 x20 0 -1
Gyc2_21 y2 0 x21 0 1
Gyc2_22 y2 0 x22 0 -1
Gyc2_23 y2 0 x23 0 1
Gyc2_24 y2 0 x24 0 0.939145106850176
Gyc2_25 y2 0 x25 0 -0.529529018022863
Gyc2_26 y2 0 x26 0 0.220740965700121
Gyc2_27 y2 0 x27 0 0.971509422487495
Gyc2_28 y2 0 x28 0 -0.0747637334494474
Gyc2_29 y2 0 x29 0 -1
Gyc2_30 y2 0 x30 0 -1
Gyc2_31 y2 0 x31 0 -1
Gyc2_32 y2 0 x32 0 0.440052770819174
Gyc2_33 y2 0 x33 0 -1
Gyc2_34 y2 0 x34 0 1
Gyc2_35 y2 0 x35 0 1
Gyc2_36 y2 0 x36 0 1
Gyc2_37 y2 0 x37 0 -1
Gyc2_38 y2 0 x38 0 1
Gyc2_39 y2 0 x39 0 -1
Gyc2_40 y2 0 x40 0 -0.947769592609844
Gyc2_41 y2 0 x41 0 -1
Gyc2_42 y2 0 x42 0 1
Gyc2_43 y2 0 x43 0 1
Gyc2_44 y2 0 x44 0 1
Gyc2_45 y2 0 x45 0 -1
Gyc2_46 y2 0 x46 0 -1
Gyc2_47 y2 0 x47 0 -1
Gyc2_48 y2 0 x48 0 -1
Gyc2_49 y2 0 x49 0 -1
Gyc2_50 y2 0 x50 0 1
Gyc2_51 y2 0 x51 0 0.513411338995705
Gyc2_52 y2 0 x52 0 -1
Gyc2_53 y2 0 x53 0 1
Gyc2_54 y2 0 x54 0 -1
Gyc2_55 y2 0 x55 0 1
Gyc2_56 y2 0 x56 0 1
Gyc2_57 y2 0 x57 0 1
Gyc2_58 y2 0 x58 0 -1
Gyc2_59 y2 0 x59 0 1
Gyc2_60 y2 0 x60 0 -1
Gyc2_61 y2 0 x61 0 1
Gyc2_62 y2 0 x62 0 -1
Gyc2_63 y2 0 x63 0 1
Gyc2_64 y2 0 x64 0 -1
Gyc2_65 y2 0 x65 0 1
Gyc2_66 y2 0 x66 0 -1
Gyc2_67 y2 0 x67 0 -1
Gyc2_68 y2 0 x68 0 1
Gyc2_69 y2 0 x69 0 -1
Gyc2_70 y2 0 x70 0 -1
Gyc2_71 y2 0 x71 0 1
Gyc2_72 y2 0 x72 0 -1
Gyc2_73 y2 0 x73 0 1
Gyc2_74 y2 0 x74 0 -1
Gyc2_75 y2 0 x75 0 1
Gyc2_76 y2 0 x76 0 1
Gyc2_77 y2 0 x77 0 1
Gyc2_78 y2 0 x78 0 -1
Gyc2_79 y2 0 x79 0 -1
Gyc2_80 y2 0 x80 0 -1
Gyc2_81 y2 0 x81 0 -1
Gyc2_82 y2 0 x82 0 -1
Gyc2_83 y2 0 x83 0 -1
Gyc2_84 y2 0 x84 0 -1
Gyc2_85 y2 0 x85 0 1
Gyc2_86 y2 0 x86 0 -1
Gyc2_87 y2 0 x87 0 1
Gyc2_88 y2 0 x88 0 -1
Gyc2_89 y2 0 x89 0 1
Gyc2_90 y2 0 x90 0 1
Gyc2_91 y2 0 x91 0 1
Gyc2_92 y2 0 x92 0 -1
Gyc2_93 y2 0 x93 0 1
Gyc2_94 y2 0 x94 0 1
Gyc2_95 y2 0 x95 0 1
Gyc2_96 y2 0 x96 0 1
Gyc2_97 y2 0 x97 0 -1
Gyc2_98 y2 0 x98 0 1
Gyc2_99 y2 0 x99 0 1
Gyc2_100 y2 0 x100 0 -1
Gyc2_101 y2 0 x101 0 1
Gyc2_102 y2 0 x102 0 1
Gyc2_103 y2 0 x103 0 -1
Gyc2_104 y2 0 x104 0 1
Gyc2_105 y2 0 x105 0 -1
Gyc2_106 y2 0 x106 0 -1
Gyc2_107 y2 0 x107 0 -1
Gyc2_108 y2 0 x108 0 1
Gyc2_109 y2 0 x109 0 1
Gyc2_110 y2 0 x110 0 1
Gyc2_111 y2 0 x111 0 1
Gyc2_112 y2 0 x112 0 1
Gyc2_113 y2 0 x113 0 -1
Gyc2_114 y2 0 x114 0 1
Gyc2_115 y2 0 x115 0 -1
Gyc2_116 y2 0 x116 0 1
Gyc2_117 y2 0 x117 0 1
Gyc2_118 y2 0 x118 0 -1
Gyc2_119 y2 0 x119 0 -1
Gyc2_120 y2 0 x120 0 1
Gyc2_121 y2 0 x121 0 1
Gyc2_122 y2 0 x122 0 -1
Gyc2_123 y2 0 x123 0 -1
Gyc2_124 y2 0 x124 0 1
Gyc2_125 y2 0 x125 0 -1
Gyc2_126 y2 0 x126 0 -1
Gyc2_127 y2 0 x127 0 -1
Gyc2_128 y2 0 x128 0 -1
Gyc2_129 y2 0 x129 0 -1
Gyc2_130 y2 0 x130 0 1
Gyc2_131 y2 0 x131 0 1
Gyc2_132 y2 0 x132 0 1
Gyc2_133 y2 0 x133 0 0.0956294252734779
Gyc2_134 y2 0 x134 0 -1
Gyc2_135 y2 0 x135 0 1
Gyc2_136 y2 0 x136 0 1
Gyc2_137 y2 0 x137 0 -1
Gyc2_138 y2 0 x138 0 1
Gyc2_139 y2 0 x139 0 1
Gyc2_140 y2 0 x140 0 -1
Gyc2_141 y2 0 x141 0 1
Gyc2_142 y2 0 x142 0 -1
Gyc2_143 y2 0 x143 0 1
Gyc2_144 y2 0 x144 0 -1
Gyc2_145 y2 0 x145 0 -1
Gyc2_146 y2 0 x146 0 1
Gyc2_147 y2 0 x147 0 -1
Gyc2_148 y2 0 x148 0 -1
Gyc2_149 y2 0 x149 0 1
Gyc2_150 y2 0 x150 0 -1
Gyc2_151 y2 0 x151 0 -1
Gyc2_152 y2 0 x152 0 1
Gyc2_153 y2 0 x153 0 1
Gyc2_154 y2 0 x154 0 1
Gyc2_155 y2 0 x155 0 1
Gyc2_156 y2 0 x156 0 1
Gyc2_157 y2 0 x157 0 1
Gyc2_158 y2 0 x158 0 -1
Gyc2_159 y2 0 x159 0 -1
Gyc2_160 y2 0 x160 0 -1
Gyc2_161 y2 0 x161 0 1
Gyc2_162 y2 0 x162 0 -1
Gyc2_163 y2 0 x163 0 -1
Gyc2_164 y2 0 x164 0 -1
Gyc2_165 y2 0 x165 0 1
Gyc2_166 y2 0 x166 0 1
Gyc2_167 y2 0 x167 0 1
Gyc2_168 y2 0 x168 0 1
Gyc2_169 y2 0 x169 0 -1
Gyc2_170 y2 0 x170 0 -1
Gyc2_171 y2 0 x171 0 1
Gyc2_172 y2 0 x172 0 1
Gyc2_173 y2 0 x173 0 -1
Gyc2_174 y2 0 x174 0 -1
Gyc2_175 y2 0 x175 0 -1
Gyc2_176 y2 0 x176 0 -1
Gyc2_177 y2 0 x177 0 -1
Gyc2_178 y2 0 x178 0 1
Gyc2_179 y2 0 x179 0 1
Gyc2_180 y2 0 x180 0 1
Gyc2_181 y2 0 x181 0 1
Gyc2_182 y2 0 x182 0 1
Gyc2_183 y2 0 x183 0 1
Gyc2_184 y2 0 x184 0 1
Gyc2_185 y2 0 x185 0 -1
Gyc2_186 y2 0 x186 0 1
Gyc2_187 y2 0 x187 0 1
Gyc2_188 y2 0 x188 0 -1
Gyc2_189 y2 0 x189 0 1
Gyc2_190 y2 0 x190 0 -1
Gyc2_191 y2 0 x191 0 1
Gyc2_192 y2 0 x192 0 -1
Gyc2_193 y2 0 x193 0 -1
Gyc2_194 y2 0 x194 0 1
Gyc2_195 y2 0 x195 0 0.148813095559048
Gyc2_196 y2 0 x196 0 1
Gyc2_197 y2 0 x197 0 -1
Gyc2_198 y2 0 x198 0 1
Gyc2_199 y2 0 x199 0 1
Gyc2_200 y2 0 x200 0 1
Gyc2_201 y2 0 x201 0 1
Gyc2_202 y2 0 x202 0 -1
Gyc2_203 y2 0 x203 0 1
Gyc2_204 y2 0 x204 0 -0.9618895514875
Gyc2_205 y2 0 x205 0 1
Gyc2_206 y2 0 x206 0 1
Gyc2_207 y2 0 x207 0 -1
Gyc2_208 y2 0 x208 0 1
Gyc2_209 y2 0 x209 0 -1
Gyc2_210 y2 0 x210 0 1
Gyc2_211 y2 0 x211 0 1
Gyc2_212 y2 0 x212 0 1
Gyc2_213 y2 0 x213 0 -1
Gyc2_214 y2 0 x214 0 1
Gyc2_215 y2 0 x215 0 -1
Gyc2_216 y2 0 x216 0 -1
Gyc2_217 y2 0 x217 0 1
Gyc2_218 y2 0 x218 0 1
Gyc2_219 y2 0 x219 0 -1
Gyc2_220 y2 0 x220 0 1
Gyc2_221 y2 0 x221 0 -1
Gyc2_222 y2 0 x222 0 0.327142461049684
Gyc2_223 y2 0 x223 0 1
Gyc2_224 y2 0 x224 0 -1
Gyc2_225 y2 0 x225 0 1
Gyc2_226 y2 0 x226 0 1
Gyc2_227 y2 0 x227 0 1
Gyc2_228 y2 0 x228 0 -1
Gyc2_229 y2 0 x229 0 1
Gyc2_230 y2 0 x230 0 1
Gyc2_231 y2 0 x231 0 -1
Gyc2_232 y2 0 x232 0 -1
Gyc2_233 y2 0 x233 0 1
Gyc2_234 y2 0 x234 0 -1
Gyc2_235 y2 0 x235 0 -1
Gyc2_236 y2 0 x236 0 -1
Gyc2_237 y2 0 x237 0 1
Gyc2_238 y2 0 x238 0 -1
Gyc2_239 y2 0 x239 0 -1
Gyc2_240 y2 0 x240 0 1
.ENDS
